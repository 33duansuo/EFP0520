`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/14 15:13:27
// Design Name: 
// Module Name: lut
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module lut_add(
    input  [4:0] m_bit1, //
    input  [4:0] m_bit2, //
    input wire [10:0]addra[3:0][7:0],
    output wire [10:0]result_bin[3:0][7:0]
    );

integer i;
integer j;
// 声明一个 wire 来存储最大位数
wire [4:0] max_bit;

// 计算 m_bit1 和 m_bit2 中的最大值
assign max_bit = (m_bit1 > m_bit2) ? m_bit1 : m_bit2;

// 声明数组
reg [31:0][4:0]M1B2;
reg [79:0][5:0]M2B2; 
reg [191:0][6:0]M3B2;
reg [447:0][7:0]M4B2;
reg [1023:0][8:0]M5B2;
reg [2303:0][9:0]M6B2;

// 声明用于存储查找结果的寄存器
reg [10:0] lookup_result_0[3:0][7:0];

initial begin
    M1B2[0] = 2;  M1B2[1] = 3;
    M1B2[2] = 2;  M1B2[3] = 3;
    M1B2[4] = 1;  M1B2[5] = 2;
    M1B2[6] = 1;  M1B2[7] = 2;
    M1B2[8] = 1;  M1B2[9] = 1;
    M1B2[10] = 1; M1B2[11] = 1;
    M1B2[12] = 0; M1B2[13] = 0;
    M1B2[14] = 0; M1B2[15] = 1;
    M1B2[16] = 12; M1B2[17] = 27;
    M1B2[18] = 12; M1B2[19] = 27;
    M1B2[20] = 28; M1B2[21] = 26;
    M1B2[22] = 28; M1B2[23] = 30;
    M1B2[24] = 29; M1B2[25] = 29;
    M1B2[26] = 29; M1B2[27] = 30;
    M1B2[28] = 30; M1B2[29] = 29;
    M1B2[30] = 30; M1B2[31] = 31;
end
initial begin
    M2B2[0] = 4;  M2B2[1] = 5;  M2B2[2] = 5;  M2B2[3] = 6;
    M2B2[4] = 4;  M2B2[5] = 5;  M2B2[6] = 5;  M2B2[7] = 6;
    M2B2[8] = 2;  M2B2[9] = 3;  M2B2[10] = 3; M2B2[11] = 4;
    M2B2[12] = 2; M2B2[13] = 3; M2B2[14] = 4; M2B2[15] = 4;
    M2B2[16] = 1; M2B2[17] = 1; M2B2[18] = 2; M2B2[19] = 2;
    M2B2[20] = 1; M2B2[21] = 2; M2B2[22] = 3; M2B2[23] = 4;
    M2B2[24] = 1; M2B2[25] = 1; M2B2[26] = 1; M2B2[27] = 1;
    M2B2[28] = 1; M2B2[29] = 2; M2B2[30] = 2; M2B2[31] = 3;
    M2B2[32] = 0; M2B2[33] = 0; M2B2[34] = 0; M2B2[35] = 1;
    M2B2[36] = 0; M2B2[37] = 1; M2B2[38] = 2; M2B2[39] = 3;
    M2B2[40] = 24; M2B2[41] = 50; M2B2[42] = 55; M2B2[43] = 58;
    M2B2[44] = 24; M2B2[45] = 50; M2B2[46] = 55; M2B2[47] = 58;
    M2B2[48] = 56; M2B2[49] = 55; M2B2[50] = 53; M2B2[51] = 49;
    M2B2[52] = 56; M2B2[53] = 58; M2B2[54] = 59; M2B2[55] = 61;
    M2B2[56] = 58; M2B2[57] = 58; M2B2[58] = 57; M2B2[59] = 57;
    M2B2[60] = 58; M2B2[61] = 60; M2B2[62] = 61; M2B2[63] = 62;
    M2B2[64] = 59; M2B2[65] = 59; M2B2[66] = 59; M2B2[67] = 59;
    M2B2[68] = 59; M2B2[69] = 60; M2B2[70] = 61; M2B2[71] = 63;
    M2B2[72] = 60; M2B2[73] = 60; M2B2[74] = 59; M2B2[75] = 59;
    M2B2[76] = 60; M2B2[77] = 61; M2B2[78] = 62; M2B2[79] = 63;
end
initial begin
    M3B2[0] = 8;   M3B2[1] = 9;   M3B2[2] = 9;   M3B2[3] = 10;
    M3B2[4] = 10;  M3B2[5] = 11;  M3B2[6] = 11;  M3B2[7] = 12;
    M3B2[8] = 8;   M3B2[9] = 9;   M3B2[10] = 9;  M3B2[11] = 10;
    M3B2[12] = 10; M3B2[13] = 11; M3B2[14] = 11; M3B2[15] = 12;
    M3B2[16] = 5;  M3B2[17] = 5;  M3B2[18] = 5;  M3B2[19] = 6;
    M3B2[20] = 6;  M3B2[21] = 7;  M3B2[22] = 7;  M3B2[23] = 8;
    M3B2[24] = 5;  M3B2[25] = 5;  M3B2[26] = 6;  M3B2[27] = 7;
    M3B2[28] = 7;  M3B2[29] = 8;  M3B2[30] = 9;  M3B2[31] = 10;
    M3B2[32] = 3;  M3B2[33] = 3;  M3B2[34] = 3;  M3B2[35] = 3;
    M3B2[36] = 3;  M3B2[37] = 4;  M3B2[38] = 4;  M3B2[39] = 4;
    M3B2[40] = 3;  M3B2[41] = 3;  M3B2[42] = 4;  M3B2[43] = 5;
    M3B2[44] = 6;  M3B2[45] = 7;  M3B2[46] = 8;  M3B2[47] = 8;
    M3B2[48] = 1;  M3B2[49] = 1;  M3B2[50] = 2;  M3B2[51] = 2;
    M3B2[52] = 2;  M3B2[53] = 2;  M3B2[54] = 2;  M3B2[55] = 2;
    M3B2[56] = 1;  M3B2[57] = 2;  M3B2[58] = 3;  M3B2[59] = 4;
    M3B2[60] = 5;  M3B2[61] = 6;  M3B2[62] = 7;  M3B2[63] = 8;
    M3B2[64] = 1;  M3B2[65] = 1;  M3B2[66] = 1;  M3B2[67] = 1;
    M3B2[68] = 1;  M3B2[69] = 1;  M3B2[70] = 1;  M3B2[71] = 1;
    M3B2[72] = 1;  M3B2[73] = 2;  M3B2[74] = 3;  M3B2[75] = 4;
    M3B2[76] = 4;  M3B2[77] = 5;  M3B2[78] = 6;  M3B2[79] = 7;
    M3B2[80] = 0;  M3B2[81] = 0;  M3B2[82] = 0;  M3B2[83] = 0;
    M3B2[84] = 0;  M3B2[85] = 1;  M3B2[86] = 1;  M3B2[87] = 1;
    M3B2[88] = 0;  M3B2[89] = 1;  M3B2[90] = 2;  M3B2[91] = 3;
    M3B2[92] = 4;  M3B2[93] = 5;  M3B2[94] = 6;  M3B2[95] = 7;
    M3B2[96] = 48;  M3B2[97] = 92;  M3B2[98] = 101; M3B2[99] = 106;
    M3B2[100] = 110; M3B2[101] = 113; M3B2[102] = 116; M3B2[103] = 118;
    M3B2[104] = 48;  M3B2[105] = 92;  M3B2[106] = 101; M3B2[107] = 106;
    M3B2[108] = 110; M3B2[109] = 113; M3B2[110] = 116; M3B2[111] = 118;
    M3B2[112] = 112; M3B2[113] = 111; M3B2[114] = 110; M3B2[115] = 108;
    M3B2[116] = 106; M3B2[117] = 103; M3B2[118] = 99;  M3B2[119] = 91;
    M3B2[120] = 112; M3B2[121] = 114; M3B2[122] = 116; M3B2[123] = 117;
    M3B2[124] = 119; M3B2[125] = 120; M3B2[126] = 122; M3B2[127] = 123;
    M3B2[128] = 117; M3B2[129] = 116; M3B2[130] = 116; M3B2[131] = 115;
    M3B2[132] = 115; M3B2[133] = 114; M3B2[134] = 114; M3B2[135] = 113;
    M3B2[136] = 117; M3B2[137] = 118; M3B2[138] = 119; M3B2[139] = 121;
    M3B2[140] = 122; M3B2[141] = 123; M3B2[142] = 124; M3B2[143] = 125;
    M3B2[144] = 118; M3B2[145] = 118; M3B2[146] = 118; M3B2[147] = 118;
    M3B2[148] = 118; M3B2[149] = 118; M3B2[150] = 117; M3B2[151] = 117;
    M3B2[152] = 118; M3B2[153] = 120; M3B2[154] = 121; M3B2[155] = 122;
    M3B2[156] = 123; M3B2[157] = 124; M3B2[158] = 125; M3B2[159] = 126;
    M3B2[160] = 119; M3B2[161] = 119; M3B2[162] = 119; M3B2[163] = 119;
    M3B2[164] = 119; M3B2[165] = 119; M3B2[166] = 119; M3B2[167] = 119;
    M3B2[168] = 119; M3B2[169] = 120; M3B2[170] = 121; M3B2[171] = 122;
    M3B2[172] = 123; M3B2[173] = 125; M3B2[174] = 126; M3B2[175] = 127;
    M3B2[176] = 120; M3B2[177] = 120; M3B2[178] = 120; M3B2[179] = 120;
    M3B2[180] = 119; M3B2[181] = 119; M3B2[182] = 119; M3B2[183] = 119;
    M3B2[184] = 120; M3B2[185] = 121; M3B2[186] = 122; M3B2[187] = 123;
    M3B2[188] = 124; M3B2[189] = 125; M3B2[190] = 126; M3B2[191] = 127;
end
initial begin
    M4B2[0] = 16;  M4B2[1] = 17;  M4B2[2] = 17;  M4B2[3] = 18;
    M4B2[4] = 18;  M4B2[5] = 19;  M4B2[6] = 19;  M4B2[7] = 20;
    M4B2[8] = 20;  M4B2[9] = 21;  M4B2[10] = 22; M4B2[11] = 22;
    M4B2[12] = 23; M4B2[13] = 23; M4B2[14] = 24; M4B2[15] = 25;
    M4B2[16] = 16; M4B2[17] = 17; M4B2[18] = 17; M4B2[19] = 18;
    M4B2[20] = 18; M4B2[21] = 19; M4B2[22] = 19; M4B2[23] = 20;
    M4B2[24] = 20; M4B2[25] = 21; M4B2[26] = 22; M4B2[27] = 22;
    M4B2[28] = 23; M4B2[29] = 23; M4B2[30] = 24; M4B2[31] = 25;
    M4B2[32] = 9;  M4B2[33] = 10; M4B2[34] = 10; M4B2[35] = 10;
    M4B2[36] = 11; M4B2[37] = 11; M4B2[38] = 12; M4B2[39] = 12;
    M4B2[40] = 12; M4B2[41] = 13; M4B2[42] = 13; M4B2[43] = 14;
    M4B2[44] = 14; M4B2[45] = 15; M4B2[46] = 15; M4B2[47] = 16;
    M4B2[48] = 9;  M4B2[49] = 10; M4B2[50] = 11; M4B2[51] = 11;
    M4B2[52] = 12; M4B2[53] = 13; M4B2[54] = 14; M4B2[55] = 14;
    M4B2[56] = 15; M4B2[57] = 16; M4B2[58] = 16; M4B2[59] = 17;
    M4B2[60] = 18; M4B2[61] = 19; M4B2[62] = 20; M4B2[63] = 20;
    M4B2[64] = 5;  M4B2[65] = 5;  M4B2[66] = 6;  M4B2[67] = 6;
    M4B2[68] = 6;  M4B2[69] = 6;  M4B2[70] = 6;  M4B2[71] = 7;
    M4B2[72] = 7;  M4B2[73] = 7;  M4B2[74] = 8;  M4B2[75] = 8;
    M4B2[76] = 8;  M4B2[77] = 8;  M4B2[78] = 9;  M4B2[79] = 9;
    M4B2[80] = 5;  M4B2[81] = 6;  M4B2[82] = 7;  M4B2[83] = 8;
    M4B2[84] = 8;  M4B2[85] = 9;  M4B2[86] = 10; M4B2[87] = 11;
    M4B2[88] = 12; M4B2[89] = 13; M4B2[90] = 13; M4B2[91] = 14;
    M4B2[92] = 15; M4B2[93] = 16; M4B2[94] = 17; M4B2[95] = 18;
    M4B2[96] = 3;  M4B2[97] = 3;  M4B2[98] = 3;  M4B2[99] = 3;
    M4B2[100] = 3; M4B2[101] = 3; M4B2[102] = 3; M4B2[103] = 4;
    M4B2[104] = 4; M4B2[105] = 4; M4B2[106] = 4; M4B2[107] = 4;
    M4B2[108] = 4; M4B2[109] = 5; M4B2[110] = 5; M4B2[111] = 5;
    M4B2[112] = 3; M4B2[113] = 4; M4B2[114] = 4; M4B2[115] = 5;
    M4B2[116] = 6; M4B2[117] = 7; M4B2[118] = 8; M4B2[119] = 9;
    M4B2[120] = 10;M4B2[121] = 11;M4B2[122] = 12;M4B2[123] = 13;
    M4B2[124] = 14;M4B2[125] = 15;M4B2[126] = 16;M4B2[127] = 16;
    M4B2[128] = 1; M4B2[129] = 1; M4B2[130] = 2; M4B2[131] = 2;
    M4B2[132] = 2; M4B2[133] = 2; M4B2[134] = 2; M4B2[135] = 2;
    M4B2[136] = 2; M4B2[137] = 2; M4B2[138] = 2; M4B2[139] = 2;
    M4B2[140] = 2; M4B2[141] = 2; M4B2[142] = 2; M4B2[143] = 3;
    M4B2[144] = 1; M4B2[145] = 2; M4B2[146] = 3; M4B2[147] = 4;
    M4B2[148] = 5; M4B2[149] = 6; M4B2[150] = 7; M4B2[151] = 8;
    M4B2[152] = 9; M4B2[153] = 10;M4B2[154] = 11;M4B2[155] = 12;
    M4B2[156] = 13;M4B2[157] = 14;M4B2[158] = 15;M4B2[159] = 16;
    M4B2[160] = 1; M4B2[161] = 1; M4B2[162] = 1; M4B2[163] = 1;
    M4B2[164] = 1; M4B2[165] = 1; M4B2[166] = 1; M4B2[167] = 1;
    M4B2[168] = 1; M4B2[169] = 1; M4B2[170] = 1; M4B2[171] = 1;
    M4B2[172] = 1; M4B2[173] = 1; M4B2[174] = 1; M4B2[175] = 1;
    M4B2[176] = 1; M4B2[177] = 2; M4B2[178] = 3; M4B2[179] = 4;
    M4B2[180] = 5; M4B2[181] = 6; M4B2[182] = 7; M4B2[183] = 8;
    M4B2[184] = 8; M4B2[185] = 9; M4B2[186] = 10;M4B2[187] = 11;
    M4B2[188] = 12;M4B2[189] = 13;M4B2[190] = 14;M4B2[191] = 15;
    M4B2[192] = 0; M4B2[193] = 0; M4B2[194] = 0; M4B2[195] = 0;
    M4B2[196] = 0; M4B2[197] = 0; M4B2[198] = 0; M4B2[199] = 0;
    M4B2[200] = 0; M4B2[201] = 1; M4B2[202] = 1; M4B2[203] = 1;
    M4B2[204] = 1; M4B2[205] = 1; M4B2[206] = 1; M4B2[207] = 1;
    M4B2[208] = 0; M4B2[209] = 1; M4B2[210] = 2; M4B2[211] = 3;
    M4B2[212] = 4; M4B2[213] = 5; M4B2[214] = 6; M4B2[215] = 7;
    M4B2[216] = 8; M4B2[217] = 9; M4B2[218] = 10;M4B2[219] = 11;
    M4B2[220] = 12;M4B2[221] = 13;M4B2[222] = 14;M4B2[223] = 15;
    M4B2[224] = 96; M4B2[225] = 168;M4B2[226] = 185;M4B2[227] = 194;
    M4B2[228] = 202;M4B2[229] = 207;M4B2[230] = 212;M4B2[231] = 216;
    M4B2[232] = 220;M4B2[233] = 223;M4B2[234] = 226;M4B2[235] = 229;
    M4B2[236] = 231;M4B2[237] = 234;M4B2[238] = 236;M4B2[239] = 238;
    M4B2[240] = 96; M4B2[241] = 168;M4B2[242] = 185;M4B2[243] = 194;
    M4B2[244] = 202;M4B2[245] = 207;M4B2[246] = 212;M4B2[247] = 216;
    M4B2[248] = 220;M4B2[249] = 223;M4B2[250] = 226;M4B2[251] = 229;
    M4B2[252] = 231;M4B2[253] = 234;M4B2[254] = 236;M4B2[255] = 238;
    M4B2[256] = 224;M4B2[257] = 223;M4B2[258] = 222;M4B2[259] = 221;
    M4B2[260] = 219;M4B2[261] = 218;M4B2[262] = 216;M4B2[263] = 214;
    M4B2[264] = 212;M4B2[265] = 209;M4B2[266] = 206;M4B2[267] = 202;
    M4B2[268] = 198;M4B2[269] = 191;M4B2[270] = 183;M4B2[271] = 167;
    M4B2[272] = 224;M4B2[273] = 226;M4B2[274] = 228;M4B2[275] = 230;
    M4B2[276] = 231;M4B2[277] = 233;M4B2[278] = 235;M4B2[279] = 236;
    M4B2[280] = 238;M4B2[281] = 239;M4B2[282] = 241;M4B2[283] = 242;
    M4B2[284] = 244;M4B2[285] = 245;M4B2[286] = 247;M4B2[287] = 248;
    M4B2[288] = 233;M4B2[289] = 233;M4B2[290] = 233;M4B2[291] = 232;
    M4B2[292] = 232;M4B2[293] = 231;M4B2[294] = 231;M4B2[295] = 230;
    M4B2[296] = 230;M4B2[297] = 229;M4B2[298] = 229;M4B2[299] = 228;
    M4B2[300] = 227;M4B2[301] = 227;M4B2[302] = 226;M4B2[303] = 225;
    M4B2[304] = 233;M4B2[305] = 235;M4B2[306] = 236;M4B2[307] = 237;
    M4B2[308] = 239;M4B2[309] = 240;M4B2[310] = 241;M4B2[311] = 242;
    M4B2[312] = 244;M4B2[313] = 245;M4B2[314] = 246;M4B2[315] = 247;
    M4B2[316] = 248;M4B2[317] = 249;M4B2[318] = 251;M4B2[319] = 252;
    M4B2[320] = 237;M4B2[321] = 237;M4B2[322] = 237;M4B2[323] = 236;
    M4B2[324] = 236;M4B2[325] = 236;M4B2[326] = 236;M4B2[327] = 236;
    M4B2[328] = 236;M4B2[329] = 235;M4B2[330] = 235;M4B2[331] = 235;
    M4B2[332] = 235;M4B2[333] = 234;M4B2[334] = 234;M4B2[335] = 234;
    M4B2[336] = 237;M4B2[337] = 238;M4B2[338] = 239;M4B2[339] = 240;
    M4B2[340] = 241;M4B2[341] = 243;M4B2[342] = 244;M4B2[343] = 245;
    M4B2[344] = 246;M4B2[345] = 247;M4B2[346] = 248;M4B2[347] = 249;
    M4B2[348] = 250;M4B2[349] = 251;M4B2[350] = 252;M4B2[351] = 253;
    M4B2[352] = 239;M4B2[353] = 238;M4B2[354] = 238;M4B2[355] = 238;
    M4B2[356] = 238;M4B2[357] = 238;M4B2[358] = 238;M4B2[359] = 238;
    M4B2[360] = 238;M4B2[361] = 238;M4B2[362] = 238;M4B2[363] = 238;
    M4B2[364] = 237;M4B2[365] = 237;M4B2[366] = 237;M4B2[367] = 237;
    M4B2[368] = 239;M4B2[369] = 240;M4B2[370] = 241;M4B2[371] = 242;
    M4B2[372] = 243;M4B2[373] = 244;M4B2[374] = 245;M4B2[375] = 246;
    M4B2[376] = 247;M4B2[377] = 248;M4B2[378] = 249;M4B2[379] = 250;
    M4B2[380] = 251;M4B2[381] = 252;M4B2[382] = 253;M4B2[383] = 254;
    M4B2[384] = 239;M4B2[385] = 239;M4B2[386] = 239;M4B2[387] = 239;
    M4B2[388] = 239;M4B2[389] = 239;M4B2[390] = 239;M4B2[391] = 239;
    M4B2[392] = 239;M4B2[393] = 239;M4B2[394] = 239;M4B2[395] = 239;
    M4B2[396] = 239;M4B2[397] = 239;M4B2[398] = 239;M4B2[399] = 239;
    M4B2[400] = 239;M4B2[401] = 240;M4B2[402] = 241;M4B2[403] = 242;
    M4B2[404] = 243;M4B2[405] = 244;M4B2[406] = 245;M4B2[407] = 246;
    M4B2[408] = 247;M4B2[409] = 249;M4B2[410] = 250;M4B2[411] = 251;
    M4B2[412] = 252;M4B2[413] = 253;M4B2[414] = 254;M4B2[415] = 255;
    M4B2[416] = 240;M4B2[417] = 240;M4B2[418] = 240;M4B2[419] = 240;
    M4B2[420] = 240;M4B2[421] = 240;M4B2[422] = 240;M4B2[423] = 240;
    M4B2[424] = 239;M4B2[425] = 239;M4B2[426] = 239;M4B2[427] = 239;
    M4B2[428] = 239;M4B2[429] = 239;M4B2[430] = 239;M4B2[431] = 239;
    M4B2[432] = 240;M4B2[433] = 241;M4B2[434] = 242;M4B2[435] = 243;
    M4B2[436] = 244;M4B2[437] = 245;M4B2[438] = 246;M4B2[439] = 247;
    M4B2[440] = 248;M4B2[441] = 249;M4B2[442] = 250;M4B2[443] = 251;
    M4B2[444] = 252;M4B2[445] = 253;M4B2[446] = 254;M4B2[447] = 255;
end
initial begin
    M5B2[0] = 32;   M5B2[1] = 33;   M5B2[2] = 33;   M5B2[3] = 34;   M5B2[4] = 34;   M5B2[5] = 35;   M5B2[6] = 35;   M5B2[7] = 36;
    M5B2[8] = 36;   M5B2[9] = 37;   M5B2[10] = 37;   M5B2[11] = 38;   M5B2[12] = 38;   M5B2[13] = 39;   M5B2[14] = 40;   M5B2[15] = 40;
    M5B2[16] = 41;   M5B2[17] = 41;   M5B2[18] = 42;   M5B2[19] = 42;   M5B2[20] = 43;   M5B2[21] = 44;   M5B2[22] = 44;   M5B2[23] = 45;
    M5B2[24] = 46;   M5B2[25] = 46;   M5B2[26] = 47;   M5B2[27] = 47;   M5B2[28] = 48;   M5B2[29] = 49;   M5B2[30] = 49;   M5B2[31] = 50;
    M5B2[32] = 32;   M5B2[33] = 33;   M5B2[34] = 33;   M5B2[35] = 34;   M5B2[36] = 34;   M5B2[37] = 35;   M5B2[38] = 35;   M5B2[39] = 36;
    M5B2[40] = 36;   M5B2[41] = 37;   M5B2[42] = 37;   M5B2[43] = 38;   M5B2[44] = 38;   M5B2[45] = 39;   M5B2[46] = 40;   M5B2[47] = 40;
    M5B2[48] = 41;   M5B2[49] = 41;   M5B2[50] = 42;   M5B2[51] = 42;   M5B2[52] = 43;   M5B2[53] = 44;   M5B2[54] = 44;   M5B2[55] = 45;
    M5B2[56] = 46;   M5B2[57] = 46;   M5B2[58] = 47;   M5B2[59] = 47;   M5B2[60] = 48;   M5B2[61] = 49;   M5B2[62] = 49;   M5B2[63] = 50;
    M5B2[64] = 19;   M5B2[65] = 19;   M5B2[66] = 19;   M5B2[67] = 20;   M5B2[68] = 20;   M5B2[69] = 20;   M5B2[70] = 21;   M5B2[71] = 21;
    M5B2[72] = 22;   M5B2[73] = 22;   M5B2[74] = 22;   M5B2[75] = 23;   M5B2[76] = 23;   M5B2[77] = 23;   M5B2[78] = 24;   M5B2[79] = 24;
    M5B2[80] = 25;   M5B2[81] = 25;   M5B2[82] = 26;   M5B2[83] = 26;   M5B2[84] = 26;   M5B2[85] = 27;   M5B2[86] = 27;   M5B2[87] = 28;
    M5B2[88] = 28;   M5B2[89] = 29;   M5B2[90] = 29;   M5B2[91] = 30;   M5B2[92] = 30;   M5B2[93] = 31;   M5B2[94] = 31;   M5B2[95] = 32;
    M5B2[96] = 19;   M5B2[97] = 19;   M5B2[98] = 20;   M5B2[99] = 21;   M5B2[100] = 21;   M5B2[101] = 22;   M5B2[102] = 23;   M5B2[103] = 23;
    M5B2[104] = 24;   M5B2[105] = 25;   M5B2[106] = 26;   M5B2[107] = 26;   M5B2[108] = 27;   M5B2[109] = 28;   M5B2[110] = 29;   M5B2[111] = 29;
    M5B2[112] = 30;   M5B2[113] = 31;   M5B2[114] = 31;   M5B2[115] = 32;   M5B2[116] = 33;   M5B2[117] = 34;   M5B2[118] = 34;   M5B2[119] = 35;
    M5B2[120] = 36;   M5B2[121] = 37;   M5B2[122] = 38;   M5B2[123] = 38;   M5B2[124] = 39;   M5B2[125] = 40;   M5B2[126] = 41;   M5B2[127] = 42;
    M5B2[128] = 10;   M5B2[129] = 11;   M5B2[130] = 11;   M5B2[131] = 11;   M5B2[132] = 11;   M5B2[133] = 11;   M5B2[134] = 12;   M5B2[135] = 12;
    M5B2[136] = 12;   M5B2[137] = 12;   M5B2[138] = 12;   M5B2[139] = 13;   M5B2[140] = 13;   M5B2[141] = 13;   M5B2[142] = 13;   M5B2[143] = 14;
    M5B2[144] = 14;   M5B2[145] = 14;   M5B2[146] = 15;   M5B2[147] = 15;   M5B2[148] = 15;   M5B2[149] = 15;   M5B2[150] = 16;   M5B2[151] = 16;
    M5B2[152] = 16;   M5B2[153] = 16;   M5B2[154] = 17;   M5B2[155] = 17;   M5B2[156] = 17;   M5B2[157] = 18;   M5B2[158] = 18;   M5B2[159] = 18;
    M5B2[160] = 10;   M5B2[161] = 11;   M5B2[162] = 12;   M5B2[163] = 13;   M5B2[164] = 14;   M5B2[165] = 14;   M5B2[166] = 15;   M5B2[167] = 16;
    M5B2[168] = 17;   M5B2[169] = 18;   M5B2[170] = 18;   M5B2[171] = 19;   M5B2[172] = 20;   M5B2[173] = 21;   M5B2[174] = 22;   M5B2[175] = 23;
    M5B2[176] = 24;   M5B2[177] = 24;   M5B2[178] = 25;   M5B2[179] = 26;   M5B2[180] = 27;   M5B2[181] = 28;   M5B2[182] = 29;   M5B2[183] = 30;
    M5B2[184] = 30;   M5B2[185] = 31;   M5B2[186] = 32;   M5B2[187] = 33;   M5B2[188] = 34;   M5B2[189] = 35;   M5B2[190] = 36;   M5B2[191] = 37;
    M5B2[192] = 5;   M5B2[193] = 6;   M5B2[194] = 6;   M5B2[195] = 6;   M5B2[196] = 6;   M5B2[197] = 6;   M5B2[198] = 6;   M5B2[199] = 6;
    M5B2[200] = 6;   M5B2[201] = 7;   M5B2[202] = 7;   M5B2[203] = 7;   M5B2[204] = 7;   M5B2[205] = 7;   M5B2[206] = 7;   M5B2[207] = 7;
    M5B2[208] = 8;   M5B2[209] = 8;   M5B2[210] = 8;   M5B2[211] = 8;   M5B2[212] = 8;   M5B2[213] = 8;   M5B2[214] = 8;   M5B2[215] = 9;
    M5B2[216] = 9;   M5B2[217] = 9;   M5B2[218] = 9;   M5B2[219] = 9;   M5B2[220] = 10;   M5B2[221] = 10;   M5B2[222] = 10;   M5B2[223] = 10;
    M5B2[224] = 5;   M5B2[225] = 6;   M5B2[226] = 7;   M5B2[227] = 8;   M5B2[228] = 9;   M5B2[229] = 10;   M5B2[230] = 11;   M5B2[231] = 12;
    M5B2[232] = 13;   M5B2[233] = 14;   M5B2[234] = 14;   M5B2[235] = 15;   M5B2[236] = 16;   M5B2[237] = 17;   M5B2[238] = 18;   M5B2[239] = 19;
    M5B2[240] = 20;   M5B2[241] = 21;   M5B2[242] = 22;   M5B2[243] = 23;   M5B2[244] = 24;   M5B2[245] = 25;   M5B2[246] = 25;   M5B2[247] = 26;
    M5B2[248] = 27;   M5B2[249] = 28;   M5B2[250] = 29;   M5B2[251] = 30;   M5B2[252] = 31;   M5B2[253] = 32;   M5B2[254] = 33;   M5B2[255] = 34;
    M5B2[256] = 3;   M5B2[257] = 3;   M5B2[258] = 3;   M5B2[259] = 3;   M5B2[260] = 3;   M5B2[261] = 3;   M5B2[262] = 3;   M5B2[263] = 3;
    M5B2[264] = 3;   M5B2[265] = 3;   M5B2[266] = 3;   M5B2[267] = 4;   M5B2[268] = 4;   M5B2[269] = 4;   M5B2[270] = 4;   M5B2[271] = 4;
    M5B2[272] = 4;   M5B2[273] = 4;   M5B2[274] = 4;   M5B2[275] = 4;   M5B2[276] = 4;   M5B2[277] = 4;   M5B2[278] = 4;   M5B2[279] = 5;
    M5B2[280] = 5;   M5B2[281] = 5;   M5B2[282] = 5;   M5B2[283] = 5;   M5B2[284] = 5;   M5B2[285] = 5;   M5B2[286] = 5;   M5B2[287] = 5;
    M5B2[288] = 3;   M5B2[289] = 4;   M5B2[290] = 5;   M5B2[291] = 6;   M5B2[292] = 7;   M5B2[293] = 8;   M5B2[294] = 8;   M5B2[295] = 9;
    M5B2[296] = 10;   M5B2[297] = 11;   M5B2[298] = 12;   M5B2[299] = 13;   M5B2[300] = 14;   M5B2[301] = 15;   M5B2[302] = 16;   M5B2[303] = 17;
    M5B2[304] = 18;   M5B2[305] = 19;   M5B2[306] = 20;   M5B2[307] = 21;   M5B2[308] = 22;   M5B2[309] = 23;   M5B2[310] = 24;   M5B2[311] = 25;
    M5B2[312] = 26;   M5B2[313] = 27;   M5B2[314] = 28;   M5B2[315] = 29;   M5B2[316] = 30;   M5B2[317] = 31;   M5B2[318] = 31;   M5B2[319] = 32;
    M5B2[320] = 1;   M5B2[321] = 1;   M5B2[322] = 1;   M5B2[323] = 2;   M5B2[324] = 2;   M5B2[325] = 2;   M5B2[326] = 2;   M5B2[327] = 2;
    M5B2[328] = 2;   M5B2[329] = 2;   M5B2[330] = 2;   M5B2[331] = 2;   M5B2[332] = 2;   M5B2[333] = 2;   M5B2[334] = 2;   M5B2[335] = 2;
    M5B2[336] = 2;   M5B2[337] = 2;   M5B2[338] = 2;   M5B2[339] = 2;   M5B2[340] = 2;   M5B2[341] = 2;   M5B2[342] = 2;   M5B2[343] = 2;
    M5B2[344] = 2;   M5B2[345] = 2;   M5B2[346] = 2;   M5B2[347] = 3;   M5B2[348] = 3;   M5B2[349] = 3;   M5B2[350] = 3;   M5B2[351] = 3;
    M5B2[352] = 1;   M5B2[353] = 2;   M5B2[354] = 3;   M5B2[355] = 4;   M5B2[356] = 5;   M5B2[357] = 6;   M5B2[358] = 7;   M5B2[359] = 8;
    M5B2[360] = 9;   M5B2[361] = 10;   M5B2[362] = 11;   M5B2[363] = 12;   M5B2[364] = 13;   M5B2[365] = 14;   M5B2[366] = 15;   M5B2[367] = 16;
    M5B2[368] = 17;   M5B2[369] = 18;   M5B2[370] = 19;   M5B2[371] = 20;   M5B2[372] = 21;   M5B2[373] = 22;   M5B2[374] = 23;   M5B2[375] = 24;
    M5B2[376] = 25;   M5B2[377] = 26;   M5B2[378] = 27;   M5B2[379] = 28;   M5B2[380] = 29;   M5B2[381] = 30;   M5B2[382] = 31;   M5B2[383] = 32;
    M5B2[384] = 1;   M5B2[385] = 1;   M5B2[386] = 1;   M5B2[387] = 1;   M5B2[388] = 1;   M5B2[389] = 1;   M5B2[390] = 1;   M5B2[391] = 1;
    M5B2[392] = 1;   M5B2[393] = 1;   M5B2[394] = 1;   M5B2[395] = 1;   M5B2[396] = 1;   M5B2[397] = 1;   M5B2[398] = 1;   M5B2[399] = 1;
    M5B2[400] = 1;   M5B2[401] = 1;   M5B2[402] = 1;   M5B2[403] = 1;   M5B2[404] = 1;   M5B2[405] = 1;   M5B2[406] = 1;   M5B2[407] = 1;
    M5B2[408] = 1;   M5B2[409] = 1;   M5B2[410] = 1;   M5B2[411] = 1;   M5B2[412] = 1;   M5B2[413] = 1;   M5B2[414] = 1;   M5B2[415] = 1;
    M5B2[416] = 1;   M5B2[417] = 2;   M5B2[418] = 3;   M5B2[419] = 4;   M5B2[420] = 5;   M5B2[421] = 6;   M5B2[422] = 7;   M5B2[423] = 8;
    M5B2[424] = 9;   M5B2[425] = 10;   M5B2[426] = 11;   M5B2[427] = 12;   M5B2[428] = 13;   M5B2[429] = 14;   M5B2[430] = 15;   M5B2[431] = 16;
    M5B2[432] = 17;   M5B2[433] = 17;   M5B2[434] = 18;   M5B2[435] = 19;   M5B2[436] = 20;   M5B2[437] = 21;   M5B2[438] = 22;   M5B2[439] = 23;
    M5B2[440] = 24;   M5B2[441] = 25;   M5B2[442] = 26;   M5B2[443] = 27;   M5B2[444] = 28;   M5B2[445] = 29;   M5B2[446] = 30;   M5B2[447] = 31;
    M5B2[448] = 0;   M5B2[449] = 0;   M5B2[450] = 0;   M5B2[451] = 0;   M5B2[452] = 0;   M5B2[453] = 0;   M5B2[454] = 0;   M5B2[455] = 0;
    M5B2[456] = 0;   M5B2[457] = 0;   M5B2[458] = 0;   M5B2[459] = 0;   M5B2[460] = 0;   M5B2[461] = 0;   M5B2[462] = 0;   M5B2[463] = 0;
    M5B2[464] = 1;   M5B2[465] = 1;   M5B2[466] = 1;   M5B2[467] = 1;   M5B2[468] = 1;   M5B2[469] = 1;   M5B2[470] = 1;   M5B2[471] = 1;
    M5B2[472] = 1;   M5B2[473] = 1;   M5B2[474] = 1;   M5B2[475] = 1;   M5B2[476] = 1;   M5B2[477] = 1;   M5B2[478] = 1;   M5B2[479] = 1;
    M5B2[480] = 0;   M5B2[481] = 1;   M5B2[482] = 2;   M5B2[483] = 3;   M5B2[484] = 4;   M5B2[485] = 5;   M5B2[486] = 6;   M5B2[487] = 7;
    M5B2[488] = 8;   M5B2[489] = 9;   M5B2[490] = 10;   M5B2[491] = 11;   M5B2[492] = 12;   M5B2[493] = 13;   M5B2[494] = 14;   M5B2[495] = 15;
    M5B2[496] = 16;   M5B2[497] = 17;   M5B2[498] = 18;   M5B2[499] = 19;   M5B2[500] = 20;   M5B2[501] = 21;   M5B2[502] = 22;   M5B2[503] = 23;
    M5B2[504] = 24;   M5B2[505] = 25;   M5B2[506] = 26;   M5B2[507] = 27;   M5B2[508] = 28;   M5B2[509] = 29;   M5B2[510] = 30;   M5B2[511] = 31;
    M5B2[512] = 192;   M5B2[513] = 304;   M5B2[514] = 336;   M5B2[515] = 355;   M5B2[516] = 369;   M5B2[517] = 380;   M5B2[518] = 389;   M5B2[519] = 396;
    M5B2[520] = 403;   M5B2[521] = 409;   M5B2[522] = 414;   M5B2[523] = 419;   M5B2[524] = 424;   M5B2[525] = 428;   M5B2[526] = 432;   M5B2[527] = 436;
    M5B2[528] = 439;   M5B2[529] = 443;   M5B2[530] = 446;   M5B2[531] = 449;   M5B2[532] = 452;   M5B2[533] = 455;   M5B2[534] = 457;   M5B2[535] = 460;
    M5B2[536] = 462;   M5B2[537] = 465;   M5B2[538] = 467;   M5B2[539] = 469;   M5B2[540] = 472;   M5B2[541] = 474;   M5B2[542] = 476;   M5B2[543] = 478;
    M5B2[544] = 192;   M5B2[545] = 304;   M5B2[546] = 336;   M5B2[547] = 355;   M5B2[548] = 369;   M5B2[549] = 380;   M5B2[550] = 389;   M5B2[551] = 396;
    M5B2[552] = 403;   M5B2[553] = 409;   M5B2[554] = 414;   M5B2[555] = 419;   M5B2[556] = 424;   M5B2[557] = 428;   M5B2[558] = 432;   M5B2[559] = 436;
    M5B2[560] = 439;   M5B2[561] = 443;   M5B2[562] = 446;   M5B2[563] = 449;   M5B2[564] = 452;   M5B2[565] = 455;   M5B2[566] = 457;   M5B2[567] = 460;
    M5B2[568] = 462;   M5B2[569] = 465;   M5B2[570] = 467;   M5B2[571] = 469;   M5B2[572] = 472;   M5B2[573] = 474;   M5B2[574] = 476;   M5B2[575] = 478;
    M5B2[576] = 448;   M5B2[577] = 447;   M5B2[578] = 446;   M5B2[579] = 445;   M5B2[580] = 444;   M5B2[581] = 442;   M5B2[582] = 441;   M5B2[583] = 440;
    M5B2[584] = 438;   M5B2[585] = 437;   M5B2[586] = 435;   M5B2[587] = 434;   M5B2[588] = 432;   M5B2[589] = 430;   M5B2[590] = 428;   M5B2[591] = 426;
    M5B2[592] = 423;   M5B2[593] = 421;   M5B2[594] = 418;   M5B2[595] = 415;   M5B2[596] = 412;   M5B2[597] = 408;   M5B2[598] = 404;   M5B2[599] = 400;
    M5B2[600] = 395;   M5B2[601] = 389;   M5B2[602] = 383;   M5B2[603] = 375;   M5B2[604] = 365;   M5B2[605] = 352;   M5B2[606] = 334;   M5B2[607] = 303;
    M5B2[608] = 448;   M5B2[609] = 450;   M5B2[610] = 452;   M5B2[611] = 454;   M5B2[612] = 456;   M5B2[613] = 458;   M5B2[614] = 459;   M5B2[615] = 461;
    M5B2[616] = 463;   M5B2[617] = 465;   M5B2[618] = 466;   M5B2[619] = 468;   M5B2[620] = 470;   M5B2[621] = 471;   M5B2[622] = 473;   M5B2[623] = 474;
    M5B2[624] = 476;   M5B2[625] = 477;   M5B2[626] = 479;   M5B2[627] = 480;   M5B2[628] = 482;   M5B2[629] = 483;   M5B2[630] = 485;   M5B2[631] = 486;
    M5B2[632] = 488;   M5B2[633] = 489;   M5B2[634] = 491;   M5B2[635] = 492;   M5B2[636] = 493;   M5B2[637] = 495;   M5B2[638] = 496;   M5B2[639] = 497;
    M5B2[640] = 467;   M5B2[641] = 466;   M5B2[642] = 466;   M5B2[643] = 466;   M5B2[644] = 465;   M5B2[645] = 465;   M5B2[646] = 465;   M5B2[647] = 464;
    M5B2[648] = 464;   M5B2[649] = 463;   M5B2[650] = 463;   M5B2[651] = 462;   M5B2[652] = 462;   M5B2[653] = 461;   M5B2[654] = 461;   M5B2[655] = 460;
    M5B2[656] = 460;   M5B2[657] = 459;   M5B2[658] = 459;   M5B2[659] = 458;   M5B2[660] = 458;   M5B2[661] = 457;   M5B2[662] = 456;   M5B2[663] = 456;
    M5B2[664] = 455;   M5B2[665] = 454;   M5B2[666] = 453;   M5B2[667] = 453;   M5B2[668] = 452;   M5B2[669] = 451;   M5B2[670] = 450;   M5B2[671] = 449;
    M5B2[672] = 467;   M5B2[673] = 468;   M5B2[674] = 469;   M5B2[675] = 471;   M5B2[676] = 472;   M5B2[677] = 473;   M5B2[678] = 475;   M5B2[679] = 476;
    M5B2[680] = 477;   M5B2[681] = 478;   M5B2[682] = 480;   M5B2[683] = 481;   M5B2[684] = 482;   M5B2[685] = 483;   M5B2[686] = 485;   M5B2[687] = 486;
    M5B2[688] = 487;   M5B2[689] = 488;   M5B2[690] = 489;   M5B2[691] = 491;   M5B2[692] = 492;   M5B2[693] = 493;   M5B2[694] = 494;   M5B2[695] = 495;
    M5B2[696] = 497;   M5B2[697] = 498;   M5B2[698] = 499;   M5B2[699] = 500;   M5B2[700] = 501;   M5B2[701] = 502;   M5B2[702] = 504;   M5B2[703] = 505;
    M5B2[704] = 474;   M5B2[705] = 474;   M5B2[706] = 474;   M5B2[707] = 473;   M5B2[708] = 473;   M5B2[709] = 473;   M5B2[710] = 473;   M5B2[711] = 473;
    M5B2[712] = 473;   M5B2[713] = 472;   M5B2[714] = 472;   M5B2[715] = 472;   M5B2[716] = 472;   M5B2[717] = 472;   M5B2[718] = 471;   M5B2[719] = 471;
    M5B2[720] = 471;   M5B2[721] = 471;   M5B2[722] = 471;   M5B2[723] = 470;   M5B2[724] = 470;   M5B2[725] = 470;   M5B2[726] = 470;   M5B2[727] = 469;
    M5B2[728] = 469;   M5B2[729] = 469;   M5B2[730] = 469;   M5B2[731] = 468;   M5B2[732] = 468;   M5B2[733] = 468;   M5B2[734] = 467;   M5B2[735] = 467;
    M5B2[736] = 474;   M5B2[737] = 475;   M5B2[738] = 476;   M5B2[739] = 477;   M5B2[740] = 478;   M5B2[741] = 480;   M5B2[742] = 481;   M5B2[743] = 482;
    M5B2[744] = 483;   M5B2[745] = 484;   M5B2[746] = 485;   M5B2[747] = 486;   M5B2[748] = 487;   M5B2[749] = 488;   M5B2[750] = 490;   M5B2[751] = 491;
    M5B2[752] = 492;   M5B2[753] = 493;   M5B2[754] = 494;   M5B2[755] = 495;   M5B2[756] = 496;   M5B2[757] = 497;   M5B2[758] = 498;   M5B2[759] = 499;
    M5B2[760] = 500;   M5B2[761] = 502;   M5B2[762] = 503;   M5B2[763] = 504;   M5B2[764] = 505;   M5B2[765] = 506;   M5B2[766] = 507;   M5B2[767] = 508;
    M5B2[768] = 477;   M5B2[769] = 477;   M5B2[770] = 477;   M5B2[771] = 477;   M5B2[772] = 477;   M5B2[773] = 477;   M5B2[774] = 477;   M5B2[775] = 477;
    M5B2[776] = 476;   M5B2[777] = 476;   M5B2[778] = 476;   M5B2[779] = 476;   M5B2[780] = 476;   M5B2[781] = 476;   M5B2[782] = 476;   M5B2[783] = 476;
    M5B2[784] = 476;   M5B2[785] = 476;   M5B2[786] = 476;   M5B2[787] = 475;   M5B2[788] = 475;   M5B2[789] = 475;   M5B2[790] = 475;   M5B2[791] = 475;
    M5B2[792] = 475;   M5B2[793] = 475;   M5B2[794] = 475;   M5B2[795] = 475;   M5B2[796] = 474;   M5B2[797] = 474;   M5B2[798] = 474;   M5B2[799] = 474;
    M5B2[800] = 477;   M5B2[801] = 478;   M5B2[802] = 479;   M5B2[803] = 480;   M5B2[804] = 481;   M5B2[805] = 482;   M5B2[806] = 483;   M5B2[807] = 484;
    M5B2[808] = 486;   M5B2[809] = 487;   M5B2[810] = 488;   M5B2[811] = 489;   M5B2[812] = 490;   M5B2[813] = 491;   M5B2[814] = 492;   M5B2[815] = 493;
    M5B2[816] = 494;   M5B2[817] = 495;   M5B2[818] = 496;   M5B2[819] = 497;   M5B2[820] = 498;   M5B2[821] = 499;   M5B2[822] = 500;   M5B2[823] = 501;
    M5B2[824] = 502;   M5B2[825] = 503;   M5B2[826] = 504;   M5B2[827] = 505;   M5B2[828] = 506;   M5B2[829] = 507;   M5B2[830] = 508;   M5B2[831] = 509;
    M5B2[832] = 479;   M5B2[833] = 478;   M5B2[834] = 478;   M5B2[835] = 478;   M5B2[836] = 478;   M5B2[837] = 478;   M5B2[838] = 478;   M5B2[839] = 478;
    M5B2[840] = 478;   M5B2[841] = 478;   M5B2[842] = 478;   M5B2[843] = 478;   M5B2[844] = 478;   M5B2[845] = 478;   M5B2[846] = 478;   M5B2[847] = 478;
    M5B2[848] = 478;   M5B2[849] = 478;   M5B2[850] = 478;   M5B2[851] = 478;   M5B2[852] = 478;   M5B2[853] = 478;   M5B2[854] = 478;   M5B2[855] = 478;
    M5B2[856] = 478;   M5B2[857] = 477;   M5B2[858] = 477;   M5B2[859] = 477;   M5B2[860] = 477;   M5B2[861] = 477;   M5B2[862] = 477;   M5B2[863] = 477;
    M5B2[864] = 479;   M5B2[865] = 480;   M5B2[866] = 481;   M5B2[867] = 482;   M5B2[868] = 483;   M5B2[869] = 484;   M5B2[870] = 485;   M5B2[871] = 486;
    M5B2[872] = 487;   M5B2[873] = 488;   M5B2[874] = 489;   M5B2[875] = 490;   M5B2[876] = 491;   M5B2[877] = 492;   M5B2[878] = 493;   M5B2[879] = 494;
    M5B2[880] = 495;   M5B2[881] = 496;   M5B2[882] = 497;   M5B2[883] = 498;   M5B2[884] = 499;   M5B2[885] = 500;   M5B2[886] = 501;   M5B2[887] = 502;
    M5B2[888] = 503;   M5B2[889] = 504;   M5B2[890] = 505;   M5B2[891] = 506;   M5B2[892] = 507;   M5B2[893] = 508;   M5B2[894] = 509;   M5B2[895] = 510;
    M5B2[896] = 479;   M5B2[897] = 479;   M5B2[898] = 479;   M5B2[899] = 479;   M5B2[900] = 479;   M5B2[901] = 479;   M5B2[902] = 479;   M5B2[903] = 479;
    M5B2[904] = 479;   M5B2[905] = 479;   M5B2[906] = 479;   M5B2[907] = 479;   M5B2[908] = 479;   M5B2[909] = 479;   M5B2[910] = 479;   M5B2[911] = 479;
    M5B2[912] = 479;   M5B2[913] = 479;   M5B2[914] = 479;   M5B2[915] = 479;   M5B2[916] = 479;   M5B2[917] = 479;   M5B2[918] = 479;   M5B2[919] = 479;
    M5B2[920] = 479;   M5B2[921] = 479;   M5B2[922] = 479;   M5B2[923] = 479;   M5B2[924] = 479;   M5B2[925] = 479;   M5B2[926] = 479;   M5B2[927] = 479;
    M5B2[928] = 479;   M5B2[929] = 480;   M5B2[930] = 481;   M5B2[931] = 482;   M5B2[932] = 483;   M5B2[933] = 484;   M5B2[934] = 485;   M5B2[935] = 486;
    M5B2[936] = 487;   M5B2[937] = 488;   M5B2[938] = 489;   M5B2[939] = 490;   M5B2[940] = 491;   M5B2[941] = 492;   M5B2[942] = 493;   M5B2[943] = 494;
    M5B2[944] = 495;   M5B2[945] = 496;   M5B2[946] = 498;   M5B2[947] = 499;   M5B2[948] = 500;   M5B2[949] = 501;   M5B2[950] = 502;   M5B2[951] = 503;
    M5B2[952] = 504;   M5B2[953] = 505;   M5B2[954] = 506;   M5B2[955] = 507;   M5B2[956] = 508;   M5B2[957] = 509;   M5B2[958] = 510;   M5B2[959] = 511;
    M5B2[960] = 480;   M5B2[961] = 480;   M5B2[962] = 480;   M5B2[963] = 480;   M5B2[964] = 480;   M5B2[965] = 480;   M5B2[966] = 480;   M5B2[967] = 480;
    M5B2[968] = 480;   M5B2[969] = 480;   M5B2[970] = 480;   M5B2[971] = 480;   M5B2[972] = 480;   M5B2[973] = 480;   M5B2[974] = 480;   M5B2[975] = 479;
    M5B2[976] = 479;   M5B2[977] = 479;   M5B2[978] = 479;   M5B2[979] = 479;   M5B2[980] = 479;   M5B2[981] = 479;   M5B2[982] = 479;   M5B2[983] = 479;
    M5B2[984] = 479;   M5B2[985] = 479;   M5B2[986] = 479;   M5B2[987] = 479;   M5B2[988] = 479;   M5B2[989] = 479;   M5B2[990] = 479;   M5B2[991] = 479;
    M5B2[992] = 480;   M5B2[993] = 481;   M5B2[994] = 482;   M5B2[995] = 483;   M5B2[996] = 484;   M5B2[997] = 485;   M5B2[998] = 486;   M5B2[999] = 487;
    M5B2[1000] = 488;   M5B2[1001] = 489;   M5B2[1002] = 490;   M5B2[1003] = 491;   M5B2[1004] = 492;   M5B2[1005] = 493;   M5B2[1006] = 494;   M5B2[1007] = 495;
    M5B2[1008] = 496;   M5B2[1009] = 497;   M5B2[1010] = 498;   M5B2[1011] = 499;   M5B2[1012] = 500;   M5B2[1013] = 501;   M5B2[1014] = 502;   M5B2[1015] = 503;
    M5B2[1016] = 504;   M5B2[1017] = 505;   M5B2[1018] = 506;   M5B2[1019] = 507;   M5B2[1020] = 508;   M5B2[1021] = 509;   M5B2[1022] = 510;   M5B2[1023] = 511;
end
initial begin
    M6B2[0] = 64;   M6B2[1] = 65;   M6B2[2] = 65;   M6B2[3] = 66;   M6B2[4] = 66;   M6B2[5] = 67;   M6B2[6] = 67;   M6B2[7] = 68;
    M6B2[8] = 68;   M6B2[9] = 69;   M6B2[10] = 69;   M6B2[11] = 70;   M6B2[12] = 70;   M6B2[13] = 71;   M6B2[14] = 71;   M6B2[15] = 72;
    M6B2[16] = 72;   M6B2[17] = 73;   M6B2[18] = 73;   M6B2[19] = 74;   M6B2[20] = 75;   M6B2[21] = 75;   M6B2[22] = 76;   M6B2[23] = 76;
    M6B2[24] = 77;   M6B2[25] = 77;   M6B2[26] = 78;   M6B2[27] = 78;   M6B2[28] = 79;   M6B2[29] = 80;   M6B2[30] = 80;   M6B2[31] = 81;
    M6B2[32] = 81;   M6B2[33] = 82;   M6B2[34] = 83;   M6B2[35] = 83;   M6B2[36] = 84;   M6B2[37] = 84;   M6B2[38] = 85;   M6B2[39] = 86;
    M6B2[40] = 86;   M6B2[41] = 87;   M6B2[42] = 87;   M6B2[43] = 88;   M6B2[44] = 89;   M6B2[45] = 89;   M6B2[46] = 90;   M6B2[47] = 90;
    M6B2[48] = 91;   M6B2[49] = 92;   M6B2[50] = 92;   M6B2[51] = 93;   M6B2[52] = 94;   M6B2[53] = 94;   M6B2[54] = 95;   M6B2[55] = 96;
    M6B2[56] = 96;   M6B2[57] = 97;   M6B2[58] = 97;   M6B2[59] = 98;   M6B2[60] = 99;   M6B2[61] = 99;   M6B2[62] = 100;   M6B2[63] = 101;
    M6B2[64] = 64;   M6B2[65] = 65;   M6B2[66] = 65;   M6B2[67] = 66;   M6B2[68] = 66;   M6B2[69] = 67;   M6B2[70] = 67;   M6B2[71] = 68;
    M6B2[72] = 68;   M6B2[73] = 69;   M6B2[74] = 69;   M6B2[75] = 70;   M6B2[76] = 70;   M6B2[77] = 71;   M6B2[78] = 71;   M6B2[79] = 72;
    M6B2[80] = 72;   M6B2[81] = 73;   M6B2[82] = 73;   M6B2[83] = 74;   M6B2[84] = 75;   M6B2[85] = 75;   M6B2[86] = 76;   M6B2[87] = 76;
    M6B2[88] = 77;   M6B2[89] = 77;   M6B2[90] = 78;   M6B2[91] = 78;   M6B2[92] = 79;   M6B2[93] = 80;   M6B2[94] = 80;   M6B2[95] = 81;
    M6B2[96] = 81;   M6B2[97] = 82;   M6B2[98] = 83;   M6B2[99] = 83;   M6B2[100] = 84;   M6B2[101] = 84;   M6B2[102] = 85;   M6B2[103] = 86;
    M6B2[104] = 86;   M6B2[105] = 87;   M6B2[106] = 87;   M6B2[107] = 88;   M6B2[108] = 89;   M6B2[109] = 89;   M6B2[110] = 90;   M6B2[111] = 90;
    M6B2[112] = 91;   M6B2[113] = 92;   M6B2[114] = 92;   M6B2[115] = 93;   M6B2[116] = 94;   M6B2[117] = 94;   M6B2[118] = 95;   M6B2[119] = 96;
    M6B2[120] = 96;   M6B2[121] = 97;   M6B2[122] = 97;   M6B2[123] = 98;   M6B2[124] = 99;   M6B2[125] = 99;   M6B2[126] = 100;   M6B2[127] = 101;
    M6B2[128] = 37;   M6B2[129] = 38;   M6B2[130] = 38;   M6B2[131] = 38;   M6B2[132] = 39;   M6B2[133] = 39;   M6B2[134] = 39;   M6B2[135] = 40;
    M6B2[136] = 40;   M6B2[137] = 41;   M6B2[138] = 41;   M6B2[139] = 41;   M6B2[140] = 42;   M6B2[141] = 42;   M6B2[142] = 42;   M6B2[143] = 43;
    M6B2[144] = 43;   M6B2[145] = 43;   M6B2[146] = 44;   M6B2[147] = 44;   M6B2[148] = 45;   M6B2[149] = 45;   M6B2[150] = 45;   M6B2[151] = 46;
    M6B2[152] = 46;   M6B2[153] = 47;   M6B2[154] = 47;   M6B2[155] = 47;   M6B2[156] = 48;   M6B2[157] = 48;   M6B2[158] = 49;   M6B2[159] = 49;
    M6B2[160] = 49;   M6B2[161] = 50;   M6B2[162] = 50;   M6B2[163] = 51;   M6B2[164] = 51;   M6B2[165] = 51;   M6B2[166] = 52;   M6B2[167] = 52;
    M6B2[168] = 53;   M6B2[169] = 53;   M6B2[170] = 54;   M6B2[171] = 54;   M6B2[172] = 55;   M6B2[173] = 55;   M6B2[174] = 55;   M6B2[175] = 56;
    M6B2[176] = 56;   M6B2[177] = 57;   M6B2[178] = 57;   M6B2[179] = 58;   M6B2[180] = 58;   M6B2[181] = 59;   M6B2[182] = 59;   M6B2[183] = 60;
    M6B2[184] = 60;   M6B2[185] = 61;   M6B2[186] = 61;   M6B2[187] = 62;   M6B2[188] = 62;   M6B2[189] = 63;   M6B2[190] = 63;   M6B2[191] = 64;
    M6B2[192] = 37;   M6B2[193] = 38;   M6B2[194] = 39;   M6B2[195] = 39;   M6B2[196] = 40;   M6B2[197] = 41;   M6B2[198] = 41;   M6B2[199] = 42;
    M6B2[200] = 43;   M6B2[201] = 44;   M6B2[202] = 44;   M6B2[203] = 45;   M6B2[204] = 46;   M6B2[205] = 46;   M6B2[206] = 47;   M6B2[207] = 48;
    M6B2[208] = 48;   M6B2[209] = 49;   M6B2[210] = 50;   M6B2[211] = 51;   M6B2[212] = 51;   M6B2[213] = 52;   M6B2[214] = 53;   M6B2[215] = 53;
    M6B2[216] = 54;   M6B2[217] = 55;   M6B2[218] = 56;   M6B2[219] = 56;   M6B2[220] = 57;   M6B2[221] = 58;   M6B2[222] = 58;   M6B2[223] = 59;
    M6B2[224] = 60;   M6B2[225] = 61;   M6B2[226] = 61;   M6B2[227] = 62;   M6B2[228] = 63;   M6B2[229] = 64;   M6B2[230] = 64;   M6B2[231] = 65;
    M6B2[232] = 66;   M6B2[233] = 67;   M6B2[234] = 67;   M6B2[235] = 68;   M6B2[236] = 69;   M6B2[237] = 70;   M6B2[238] = 70;   M6B2[239] = 71;
    M6B2[240] = 72;   M6B2[241] = 73;   M6B2[242] = 74;   M6B2[243] = 74;   M6B2[244] = 75;   M6B2[245] = 76;   M6B2[246] = 77;   M6B2[247] = 77;
    M6B2[248] = 78;   M6B2[249] = 79;   M6B2[250] = 80;   M6B2[251] = 81;   M6B2[252] = 81;   M6B2[253] = 82;   M6B2[254] = 83;   M6B2[255] = 84;
    M6B2[256] = 21;   M6B2[257] = 21;   M6B2[258] = 21;   M6B2[259] = 21;   M6B2[260] = 21;   M6B2[261] = 22;   M6B2[262] = 22;   M6B2[263] = 22;
    M6B2[264] = 22;   M6B2[265] = 22;   M6B2[266] = 23;   M6B2[267] = 23;   M6B2[268] = 23;   M6B2[269] = 23;   M6B2[270] = 24;   M6B2[271] = 24;
    M6B2[272] = 24;   M6B2[273] = 24;   M6B2[274] = 24;   M6B2[275] = 25;   M6B2[276] = 25;   M6B2[277] = 25;   M6B2[278] = 25;   M6B2[279] = 26;
    M6B2[280] = 26;   M6B2[281] = 26;   M6B2[282] = 26;   M6B2[283] = 27;   M6B2[284] = 27;   M6B2[285] = 27;   M6B2[286] = 27;   M6B2[287] = 28;
    M6B2[288] = 28;   M6B2[289] = 28;   M6B2[290] = 28;   M6B2[291] = 29;   M6B2[292] = 29;   M6B2[293] = 29;   M6B2[294] = 30;   M6B2[295] = 30;
    M6B2[296] = 30;   M6B2[297] = 30;   M6B2[298] = 31;   M6B2[299] = 31;   M6B2[300] = 31;   M6B2[301] = 32;   M6B2[302] = 32;   M6B2[303] = 32;
    M6B2[304] = 32;   M6B2[305] = 33;   M6B2[306] = 33;   M6B2[307] = 33;   M6B2[308] = 34;   M6B2[309] = 34;   M6B2[310] = 34;   M6B2[311] = 35;
    M6B2[312] = 35;   M6B2[313] = 35;   M6B2[314] = 35;   M6B2[315] = 36;   M6B2[316] = 36;   M6B2[317] = 36;   M6B2[318] = 37;   M6B2[319] = 37;
    M6B2[320] = 21;   M6B2[321] = 21;   M6B2[322] = 22;   M6B2[323] = 23;   M6B2[324] = 24;   M6B2[325] = 25;   M6B2[326] = 25;   M6B2[327] = 26;
    M6B2[328] = 27;   M6B2[329] = 28;   M6B2[330] = 29;   M6B2[331] = 30;   M6B2[332] = 30;   M6B2[333] = 31;   M6B2[334] = 32;   M6B2[335] = 33;
    M6B2[336] = 34;   M6B2[337] = 34;   M6B2[338] = 35;   M6B2[339] = 36;   M6B2[340] = 37;   M6B2[341] = 38;   M6B2[342] = 39;   M6B2[343] = 39;
    M6B2[344] = 40;   M6B2[345] = 41;   M6B2[346] = 42;   M6B2[347] = 43;   M6B2[348] = 44;   M6B2[349] = 44;   M6B2[350] = 45;   M6B2[351] = 46;
    M6B2[352] = 47;   M6B2[353] = 48;   M6B2[354] = 49;   M6B2[355] = 50;   M6B2[356] = 50;   M6B2[357] = 51;   M6B2[358] = 52;   M6B2[359] = 53;
    M6B2[360] = 54;   M6B2[361] = 55;   M6B2[362] = 56;   M6B2[363] = 56;   M6B2[364] = 57;   M6B2[365] = 58;   M6B2[366] = 59;   M6B2[367] = 60;
    M6B2[368] = 61;   M6B2[369] = 62;   M6B2[370] = 63;   M6B2[371] = 63;   M6B2[372] = 64;   M6B2[373] = 65;   M6B2[374] = 66;   M6B2[375] = 67;
    M6B2[376] = 68;   M6B2[377] = 69;   M6B2[378] = 70;   M6B2[379] = 70;   M6B2[380] = 71;   M6B2[381] = 72;   M6B2[382] = 73;   M6B2[383] = 74;
    M6B2[384] = 11;   M6B2[385] = 11;   M6B2[386] = 11;   M6B2[387] = 11;   M6B2[388] = 11;   M6B2[389] = 11;   M6B2[390] = 12;   M6B2[391] = 12;
    M6B2[392] = 12;   M6B2[393] = 12;   M6B2[394] = 12;   M6B2[395] = 12;   M6B2[396] = 12;   M6B2[397] = 12;   M6B2[398] = 13;   M6B2[399] = 13;
    M6B2[400] = 13;   M6B2[401] = 13;   M6B2[402] = 13;   M6B2[403] = 13;   M6B2[404] = 13;   M6B2[405] = 13;   M6B2[406] = 14;   M6B2[407] = 14;
    M6B2[408] = 14;   M6B2[409] = 14;   M6B2[410] = 14;   M6B2[411] = 14;   M6B2[412] = 14;   M6B2[413] = 15;   M6B2[414] = 15;   M6B2[415] = 15;
    M6B2[416] = 15;   M6B2[417] = 15;   M6B2[418] = 15;   M6B2[419] = 15;   M6B2[420] = 16;   M6B2[421] = 16;   M6B2[422] = 16;   M6B2[423] = 16;
    M6B2[424] = 16;   M6B2[425] = 16;   M6B2[426] = 17;   M6B2[427] = 17;   M6B2[428] = 17;   M6B2[429] = 17;   M6B2[430] = 17;   M6B2[431] = 17;
    M6B2[432] = 18;   M6B2[433] = 18;   M6B2[434] = 18;   M6B2[435] = 18;   M6B2[436] = 18;   M6B2[437] = 19;   M6B2[438] = 19;   M6B2[439] = 19;
    M6B2[440] = 19;   M6B2[441] = 19;   M6B2[442] = 19;   M6B2[443] = 20;   M6B2[444] = 20;   M6B2[445] = 20;   M6B2[446] = 20;   M6B2[447] = 20;
    M6B2[448] = 11;   M6B2[449] = 12;   M6B2[450] = 13;   M6B2[451] = 14;   M6B2[452] = 14;   M6B2[453] = 15;   M6B2[454] = 16;   M6B2[455] = 17;
    M6B2[456] = 18;   M6B2[457] = 19;   M6B2[458] = 20;   M6B2[459] = 21;   M6B2[460] = 22;   M6B2[461] = 23;   M6B2[462] = 23;   M6B2[463] = 24;
    M6B2[464] = 25;   M6B2[465] = 26;   M6B2[466] = 27;   M6B2[467] = 28;   M6B2[468] = 29;   M6B2[469] = 30;   M6B2[470] = 31;   M6B2[471] = 32;
    M6B2[472] = 32;   M6B2[473] = 33;   M6B2[474] = 34;   M6B2[475] = 35;   M6B2[476] = 36;   M6B2[477] = 37;   M6B2[478] = 38;   M6B2[479] = 39;
    M6B2[480] = 40;   M6B2[481] = 41;   M6B2[482] = 42;   M6B2[483] = 43;   M6B2[484] = 44;   M6B2[485] = 44;   M6B2[486] = 45;   M6B2[487] = 46;
    M6B2[488] = 47;   M6B2[489] = 48;   M6B2[490] = 49;   M6B2[491] = 50;   M6B2[492] = 51;   M6B2[493] = 52;   M6B2[494] = 53;   M6B2[495] = 54;
    M6B2[496] = 55;   M6B2[497] = 56;   M6B2[498] = 56;   M6B2[499] = 57;   M6B2[500] = 58;   M6B2[501] = 59;   M6B2[502] = 60;   M6B2[503] = 61;
    M6B2[504] = 62;   M6B2[505] = 63;   M6B2[506] = 64;   M6B2[507] = 65;   M6B2[508] = 66;   M6B2[509] = 67;   M6B2[510] = 68;   M6B2[511] = 69;
    M6B2[512] = 6;   M6B2[513] = 6;   M6B2[514] = 6;   M6B2[515] = 6;   M6B2[516] = 6;   M6B2[517] = 6;   M6B2[518] = 6;   M6B2[519] = 6;
    M6B2[520] = 6;   M6B2[521] = 6;   M6B2[522] = 6;   M6B2[523] = 6;   M6B2[524] = 6;   M6B2[525] = 6;   M6B2[526] = 6;   M6B2[527] = 7;
    M6B2[528] = 7;   M6B2[529] = 7;   M6B2[530] = 7;   M6B2[531] = 7;   M6B2[532] = 7;   M6B2[533] = 7;   M6B2[534] = 7;   M6B2[535] = 7;
    M6B2[536] = 7;   M6B2[537] = 7;   M6B2[538] = 7;   M6B2[539] = 7;   M6B2[540] = 8;   M6B2[541] = 8;   M6B2[542] = 8;   M6B2[543] = 8;
    M6B2[544] = 8;   M6B2[545] = 8;   M6B2[546] = 8;   M6B2[547] = 8;   M6B2[548] = 8;   M6B2[549] = 8;   M6B2[550] = 8;   M6B2[551] = 8;
    M6B2[552] = 8;   M6B2[553] = 9;   M6B2[554] = 9;   M6B2[555] = 9;   M6B2[556] = 9;   M6B2[557] = 9;   M6B2[558] = 9;   M6B2[559] = 9;
    M6B2[560] = 9;   M6B2[561] = 9;   M6B2[562] = 9;   M6B2[563] = 10;   M6B2[564] = 10;   M6B2[565] = 10;   M6B2[566] = 10;   M6B2[567] = 10;
    M6B2[568] = 10;   M6B2[569] = 10;   M6B2[570] = 10;   M6B2[571] = 10;   M6B2[572] = 10;   M6B2[573] = 11;   M6B2[574] = 11;   M6B2[575] = 11;
    M6B2[576] = 6;   M6B2[577] = 7;   M6B2[578] = 7;   M6B2[579] = 8;   M6B2[580] = 9;   M6B2[581] = 10;   M6B2[582] = 11;   M6B2[583] = 12;
    M6B2[584] = 13;   M6B2[585] = 14;   M6B2[586] = 15;   M6B2[587] = 16;   M6B2[588] = 17;   M6B2[589] = 18;   M6B2[590] = 19;   M6B2[591] = 20;
    M6B2[592] = 21;   M6B2[593] = 22;   M6B2[594] = 23;   M6B2[595] = 24;   M6B2[596] = 25;   M6B2[597] = 25;   M6B2[598] = 26;   M6B2[599] = 27;
    M6B2[600] = 28;   M6B2[601] = 29;   M6B2[602] = 30;   M6B2[603] = 31;   M6B2[604] = 32;   M6B2[605] = 33;   M6B2[606] = 34;   M6B2[607] = 35;
    M6B2[608] = 36;   M6B2[609] = 37;   M6B2[610] = 38;   M6B2[611] = 39;   M6B2[612] = 40;   M6B2[613] = 41;   M6B2[614] = 42;   M6B2[615] = 43;
    M6B2[616] = 44;   M6B2[617] = 45;   M6B2[618] = 46;   M6B2[619] = 47;   M6B2[620] = 48;   M6B2[621] = 48;   M6B2[622] = 49;   M6B2[623] = 50;
    M6B2[624] = 51;   M6B2[625] = 52;   M6B2[626] = 53;   M6B2[627] = 54;   M6B2[628] = 55;   M6B2[629] = 56;   M6B2[630] = 57;   M6B2[631] = 58;
    M6B2[632] = 59;   M6B2[633] = 60;   M6B2[634] = 61;   M6B2[635] = 62;   M6B2[636] = 63;   M6B2[637] = 64;   M6B2[638] = 65;   M6B2[639] = 66;
    M6B2[640] = 3;   M6B2[641] = 3;   M6B2[642] = 3;   M6B2[643] = 3;   M6B2[644] = 3;   M6B2[645] = 3;   M6B2[646] = 3;   M6B2[647] = 3;
    M6B2[648] = 3;   M6B2[649] = 3;   M6B2[650] = 3;   M6B2[651] = 3;   M6B2[652] = 3;   M6B2[653] = 3;   M6B2[654] = 3;   M6B2[655] = 3;
    M6B2[656] = 3;   M6B2[657] = 3;   M6B2[658] = 3;   M6B2[659] = 3;   M6B2[660] = 4;   M6B2[661] = 4;   M6B2[662] = 4;   M6B2[663] = 4;
    M6B2[664] = 4;   M6B2[665] = 4;   M6B2[666] = 4;   M6B2[667] = 4;   M6B2[668] = 4;   M6B2[669] = 4;   M6B2[670] = 4;   M6B2[671] = 4;
    M6B2[672] = 4;   M6B2[673] = 4;   M6B2[674] = 4;   M6B2[675] = 4;   M6B2[676] = 4;   M6B2[677] = 4;   M6B2[678] = 4;   M6B2[679] = 4;
    M6B2[680] = 4;   M6B2[681] = 4;   M6B2[682] = 4;   M6B2[683] = 4;   M6B2[684] = 5;   M6B2[685] = 5;   M6B2[686] = 5;   M6B2[687] = 5;
    M6B2[688] = 5;   M6B2[689] = 5;   M6B2[690] = 5;   M6B2[691] = 5;   M6B2[692] = 5;   M6B2[693] = 5;   M6B2[694] = 5;   M6B2[695] = 5;
    M6B2[696] = 5;   M6B2[697] = 5;   M6B2[698] = 5;   M6B2[699] = 5;   M6B2[700] = 5;   M6B2[701] = 5;   M6B2[702] = 5;   M6B2[703] = 6;
    M6B2[704] = 3;   M6B2[705] = 4;   M6B2[706] = 5;   M6B2[707] = 6;   M6B2[708] = 7;   M6B2[709] = 8;   M6B2[710] = 9;   M6B2[711] = 10;
    M6B2[712] = 11;   M6B2[713] = 12;   M6B2[714] = 13;   M6B2[715] = 14;   M6B2[716] = 14;   M6B2[717] = 15;   M6B2[718] = 16;   M6B2[719] = 17;
    M6B2[720] = 18;   M6B2[721] = 19;   M6B2[722] = 20;   M6B2[723] = 21;   M6B2[724] = 22;   M6B2[725] = 23;   M6B2[726] = 24;   M6B2[727] = 25;
    M6B2[728] = 26;   M6B2[729] = 27;   M6B2[730] = 28;   M6B2[731] = 29;   M6B2[732] = 30;   M6B2[733] = 31;   M6B2[734] = 32;   M6B2[735] = 33;
    M6B2[736] = 34;   M6B2[737] = 35;   M6B2[738] = 36;   M6B2[739] = 37;   M6B2[740] = 38;   M6B2[741] = 39;   M6B2[742] = 40;   M6B2[743] = 41;
    M6B2[744] = 42;   M6B2[745] = 43;   M6B2[746] = 44;   M6B2[747] = 45;   M6B2[748] = 46;   M6B2[749] = 47;   M6B2[750] = 48;   M6B2[751] = 49;
    M6B2[752] = 50;   M6B2[753] = 51;   M6B2[754] = 52;   M6B2[755] = 53;   M6B2[756] = 54;   M6B2[757] = 55;   M6B2[758] = 56;   M6B2[759] = 57;
    M6B2[760] = 58;   M6B2[761] = 59;   M6B2[762] = 60;   M6B2[763] = 61;   M6B2[764] = 61;   M6B2[765] = 62;   M6B2[766] = 63;   M6B2[767] = 64;
    M6B2[768] = 1;   M6B2[769] = 1;   M6B2[770] = 1;   M6B2[771] = 1;   M6B2[772] = 1;   M6B2[773] = 2;   M6B2[774] = 2;   M6B2[775] = 2;
    M6B2[776] = 2;   M6B2[777] = 2;   M6B2[778] = 2;   M6B2[779] = 2;   M6B2[780] = 2;   M6B2[781] = 2;   M6B2[782] = 2;   M6B2[783] = 2;
    M6B2[784] = 2;   M6B2[785] = 2;   M6B2[786] = 2;   M6B2[787] = 2;   M6B2[788] = 2;   M6B2[789] = 2;   M6B2[790] = 2;   M6B2[791] = 2;
    M6B2[792] = 2;   M6B2[793] = 2;   M6B2[794] = 2;   M6B2[795] = 2;   M6B2[796] = 2;   M6B2[797] = 2;   M6B2[798] = 2;   M6B2[799] = 2;
    M6B2[800] = 2;   M6B2[801] = 2;   M6B2[802] = 2;   M6B2[803] = 2;   M6B2[804] = 2;   M6B2[805] = 2;   M6B2[806] = 2;   M6B2[807] = 2;
    M6B2[808] = 2;   M6B2[809] = 2;   M6B2[810] = 2;   M6B2[811] = 2;   M6B2[812] = 2;   M6B2[813] = 2;   M6B2[814] = 2;   M6B2[815] = 2;
    M6B2[816] = 2;   M6B2[817] = 2;   M6B2[818] = 2;   M6B2[819] = 2;   M6B2[820] = 2;   M6B2[821] = 3;   M6B2[822] = 3;   M6B2[823] = 3;
    M6B2[824] = 3;   M6B2[825] = 3;   M6B2[826] = 3;   M6B2[827] = 3;   M6B2[828] = 3;   M6B2[829] = 3;   M6B2[830] = 3;   M6B2[831] = 3;
    M6B2[832] = 1;   M6B2[833] = 2;   M6B2[834] = 3;   M6B2[835] = 4;   M6B2[836] = 5;   M6B2[837] = 6;   M6B2[838] = 7;   M6B2[839] = 8;
    M6B2[840] = 9;   M6B2[841] = 10;   M6B2[842] = 11;   M6B2[843] = 12;   M6B2[844] = 13;   M6B2[845] = 14;   M6B2[846] = 15;   M6B2[847] = 16;
    M6B2[848] = 17;   M6B2[849] = 18;   M6B2[850] = 19;   M6B2[851] = 20;   M6B2[852] = 21;   M6B2[853] = 22;   M6B2[854] = 23;   M6B2[855] = 24;
    M6B2[856] = 25;   M6B2[857] = 26;   M6B2[858] = 27;   M6B2[859] = 28;   M6B2[860] = 29;   M6B2[861] = 30;   M6B2[862] = 31;   M6B2[863] = 32;
    M6B2[864] = 33;   M6B2[865] = 34;   M6B2[866] = 35;   M6B2[867] = 36;   M6B2[868] = 37;   M6B2[869] = 38;   M6B2[870] = 39;   M6B2[871] = 40;
    M6B2[872] = 41;   M6B2[873] = 42;   M6B2[874] = 43;   M6B2[875] = 44;   M6B2[876] = 45;   M6B2[877] = 46;   M6B2[878] = 47;   M6B2[879] = 48;
    M6B2[880] = 49;   M6B2[881] = 50;   M6B2[882] = 51;   M6B2[883] = 52;   M6B2[884] = 53;   M6B2[885] = 54;   M6B2[886] = 55;   M6B2[887] = 56;
    M6B2[888] = 57;   M6B2[889] = 58;   M6B2[890] = 59;   M6B2[891] = 60;   M6B2[892] = 61;   M6B2[893] = 62;   M6B2[894] = 63;   M6B2[895] = 64;
    M6B2[896] = 1;   M6B2[897] = 1;   M6B2[898] = 1;   M6B2[899] = 1;   M6B2[900] = 1;   M6B2[901] = 1;   M6B2[902] = 1;   M6B2[903] = 1;
    M6B2[904] = 1;   M6B2[905] = 1;   M6B2[906] = 1;   M6B2[907] = 1;   M6B2[908] = 1;   M6B2[909] = 1;   M6B2[910] = 1;   M6B2[911] = 1;
    M6B2[912] = 1;   M6B2[913] = 1;   M6B2[914] = 1;   M6B2[915] = 1;   M6B2[916] = 1;   M6B2[917] = 1;   M6B2[918] = 1;   M6B2[919] = 1;
    M6B2[920] = 1;   M6B2[921] = 1;   M6B2[922] = 1;   M6B2[923] = 1;   M6B2[924] = 1;   M6B2[925] = 1;   M6B2[926] = 1;   M6B2[927] = 1;
    M6B2[928] = 1;   M6B2[929] = 1;   M6B2[930] = 1;   M6B2[931] = 1;   M6B2[932] = 1;   M6B2[933] = 1;   M6B2[934] = 1;   M6B2[935] = 1;
    M6B2[936] = 1;   M6B2[937] = 1;   M6B2[938] = 1;   M6B2[939] = 1;   M6B2[940] = 1;   M6B2[941] = 1;   M6B2[942] = 1;   M6B2[943] = 1;
    M6B2[944] = 1;   M6B2[945] = 1;   M6B2[946] = 1;   M6B2[947] = 1;   M6B2[948] = 1;   M6B2[949] = 1;   M6B2[950] = 1;   M6B2[951] = 1;
    M6B2[952] = 1;   M6B2[953] = 1;   M6B2[954] = 1;   M6B2[955] = 1;   M6B2[956] = 1;   M6B2[957] = 1;   M6B2[958] = 1;   M6B2[959] = 1;
    M6B2[960] = 1;   M6B2[961] = 2;   M6B2[962] = 3;   M6B2[963] = 4;   M6B2[964] = 5;   M6B2[965] = 6;   M6B2[966] = 7;   M6B2[967] = 8;
    M6B2[968] = 9;   M6B2[969] = 10;   M6B2[970] = 11;   M6B2[971] = 12;   M6B2[972] = 13;   M6B2[973] = 14;   M6B2[974] = 15;   M6B2[975] = 16;
    M6B2[976] = 17;   M6B2[977] = 18;   M6B2[978] = 19;   M6B2[979] = 20;   M6B2[980] = 21;   M6B2[981] = 22;   M6B2[982] = 23;   M6B2[983] = 24;
    M6B2[984] = 25;   M6B2[985] = 26;   M6B2[986] = 27;   M6B2[987] = 28;   M6B2[988] = 29;   M6B2[989] = 30;   M6B2[990] = 31;   M6B2[991] = 32;
    M6B2[992] = 33;   M6B2[993] = 34;   M6B2[994] = 34;   M6B2[995] = 35;   M6B2[996] = 36;   M6B2[997] = 37;   M6B2[998] = 38;   M6B2[999] = 39;
    M6B2[1000] = 40;   M6B2[1001] = 41;   M6B2[1002] = 42;   M6B2[1003] = 43;   M6B2[1004] = 44;   M6B2[1005] = 45;   M6B2[1006] = 46;   M6B2[1007] = 47;
    M6B2[1008] = 48;   M6B2[1009] = 49;   M6B2[1010] = 50;   M6B2[1011] = 51;   M6B2[1012] = 52;   M6B2[1013] = 53;   M6B2[1014] = 54;   M6B2[1015] = 55;
    M6B2[1016] = 56;   M6B2[1017] = 57;   M6B2[1018] = 58;   M6B2[1019] = 59;   M6B2[1020] = 60;   M6B2[1021] = 61;   M6B2[1022] = 62;   M6B2[1023] = 63;
    M6B2[1024] = 0;   M6B2[1025] = 0;   M6B2[1026] = 0;   M6B2[1027] = 0;   M6B2[1028] = 0;   M6B2[1029] = 0;   M6B2[1030] = 0;   M6B2[1031] = 0;
    M6B2[1032] = 0;   M6B2[1033] = 0;   M6B2[1034] = 0;   M6B2[1035] = 0;   M6B2[1036] = 0;   M6B2[1037] = 0;   M6B2[1038] = 0;   M6B2[1039] = 0;
    M6B2[1040] = 0;   M6B2[1041] = 0;   M6B2[1042] = 0;   M6B2[1043] = 0;   M6B2[1044] = 0;   M6B2[1045] = 0;   M6B2[1046] = 0;   M6B2[1047] = 0;
    M6B2[1048] = 0;   M6B2[1049] = 0;   M6B2[1050] = 0;   M6B2[1051] = 0;   M6B2[1052] = 0;   M6B2[1053] = 0;   M6B2[1054] = 0;   M6B2[1055] = 1;
    M6B2[1056] = 1;   M6B2[1057] = 1;   M6B2[1058] = 1;   M6B2[1059] = 1;   M6B2[1060] = 1;   M6B2[1061] = 1;   M6B2[1062] = 1;   M6B2[1063] = 1;
    M6B2[1064] = 1;   M6B2[1065] = 1;   M6B2[1066] = 1;   M6B2[1067] = 1;   M6B2[1068] = 1;   M6B2[1069] = 1;   M6B2[1070] = 1;   M6B2[1071] = 1;
    M6B2[1072] = 1;   M6B2[1073] = 1;   M6B2[1074] = 1;   M6B2[1075] = 1;   M6B2[1076] = 1;   M6B2[1077] = 1;   M6B2[1078] = 1;   M6B2[1079] = 1;
    M6B2[1080] = 1;   M6B2[1081] = 1;   M6B2[1082] = 1;   M6B2[1083] = 1;   M6B2[1084] = 1;   M6B2[1085] = 1;   M6B2[1086] = 1;   M6B2[1087] = 1;
    M6B2[1088] = 0;   M6B2[1089] = 1;   M6B2[1090] = 2;   M6B2[1091] = 3;   M6B2[1092] = 4;   M6B2[1093] = 5;   M6B2[1094] = 6;   M6B2[1095] = 7;
    M6B2[1096] = 8;   M6B2[1097] = 9;   M6B2[1098] = 10;   M6B2[1099] = 11;   M6B2[1100] = 12;   M6B2[1101] = 13;   M6B2[1102] = 14;   M6B2[1103] = 15;
    M6B2[1104] = 16;   M6B2[1105] = 17;   M6B2[1106] = 18;   M6B2[1107] = 19;   M6B2[1108] = 20;   M6B2[1109] = 21;   M6B2[1110] = 22;   M6B2[1111] = 23;
    M6B2[1112] = 24;   M6B2[1113] = 25;   M6B2[1114] = 26;   M6B2[1115] = 27;   M6B2[1116] = 28;   M6B2[1117] = 29;   M6B2[1118] = 30;   M6B2[1119] = 31;
    M6B2[1120] = 32;   M6B2[1121] = 33;   M6B2[1122] = 34;   M6B2[1123] = 35;   M6B2[1124] = 36;   M6B2[1125] = 37;   M6B2[1126] = 38;   M6B2[1127] = 39;
    M6B2[1128] = 40;   M6B2[1129] = 41;   M6B2[1130] = 42;   M6B2[1131] = 43;   M6B2[1132] = 44;   M6B2[1133] = 45;   M6B2[1134] = 46;   M6B2[1135] = 47;
    M6B2[1136] = 48;   M6B2[1137] = 49;   M6B2[1138] = 50;   M6B2[1139] = 51;   M6B2[1140] = 52;   M6B2[1141] = 53;   M6B2[1142] = 54;   M6B2[1143] = 55;
    M6B2[1144] = 56;   M6B2[1145] = 57;   M6B2[1146] = 58;   M6B2[1147] = 59;   M6B2[1148] = 60;   M6B2[1149] = 61;   M6B2[1150] = 62;   M6B2[1151] = 63;
    M6B2[1152] = 384;   M6B2[1153] = 543;   M6B2[1154] = 607;   M6B2[1155] = 645;   M6B2[1156] = 672;   M6B2[1157] = 693;   M6B2[1158] = 711;   M6B2[1159] = 725;
    M6B2[1160] = 738;   M6B2[1161] = 750;   M6B2[1162] = 760;   M6B2[1163] = 769;   M6B2[1164] = 778;   M6B2[1165] = 786;   M6B2[1166] = 793;   M6B2[1167] = 800;
    M6B2[1168] = 806;   M6B2[1169] = 812;   M6B2[1170] = 818;   M6B2[1171] = 824;   M6B2[1172] = 829;   M6B2[1173] = 834;   M6B2[1174] = 839;   M6B2[1175] = 843;
    M6B2[1176] = 848;   M6B2[1177] = 852;   M6B2[1178] = 856;   M6B2[1179] = 860;   M6B2[1180] = 864;   M6B2[1181] = 868;   M6B2[1182] = 872;   M6B2[1183] = 875;
    M6B2[1184] = 879;   M6B2[1185] = 882;   M6B2[1186] = 885;   M6B2[1187] = 888;   M6B2[1188] = 892;   M6B2[1189] = 895;   M6B2[1190] = 898;   M6B2[1191] = 901;
    M6B2[1192] = 903;   M6B2[1193] = 906;   M6B2[1194] = 909;   M6B2[1195] = 912;   M6B2[1196] = 914;   M6B2[1197] = 917;   M6B2[1198] = 920;   M6B2[1199] = 922;
    M6B2[1200] = 925;   M6B2[1201] = 927;   M6B2[1202] = 929;   M6B2[1203] = 932;   M6B2[1204] = 934;   M6B2[1205] = 937;   M6B2[1206] = 939;   M6B2[1207] = 941;
    M6B2[1208] = 943;   M6B2[1209] = 945;   M6B2[1210] = 948;   M6B2[1211] = 950;   M6B2[1212] = 952;   M6B2[1213] = 954;   M6B2[1214] = 956;   M6B2[1215] = 958;
    M6B2[1216] = 384;   M6B2[1217] = 543;   M6B2[1218] = 607;   M6B2[1219] = 645;   M6B2[1220] = 672;   M6B2[1221] = 693;   M6B2[1222] = 711;   M6B2[1223] = 725;
    M6B2[1224] = 738;   M6B2[1225] = 750;   M6B2[1226] = 760;   M6B2[1227] = 769;   M6B2[1228] = 778;   M6B2[1229] = 786;   M6B2[1230] = 793;   M6B2[1231] = 800;
    M6B2[1232] = 806;   M6B2[1233] = 812;   M6B2[1234] = 818;   M6B2[1235] = 824;   M6B2[1236] = 829;   M6B2[1237] = 834;   M6B2[1238] = 839;   M6B2[1239] = 843;
    M6B2[1240] = 848;   M6B2[1241] = 852;   M6B2[1242] = 856;   M6B2[1243] = 860;   M6B2[1244] = 864;   M6B2[1245] = 868;   M6B2[1246] = 872;   M6B2[1247] = 875;
    M6B2[1248] = 879;   M6B2[1249] = 882;   M6B2[1250] = 885;   M6B2[1251] = 888;   M6B2[1252] = 892;   M6B2[1253] = 895;   M6B2[1254] = 898;   M6B2[1255] = 901;
    M6B2[1256] = 903;   M6B2[1257] = 906;   M6B2[1258] = 909;   M6B2[1259] = 912;   M6B2[1260] = 914;   M6B2[1261] = 917;   M6B2[1262] = 920;   M6B2[1263] = 922;
    M6B2[1264] = 925;   M6B2[1265] = 927;   M6B2[1266] = 929;   M6B2[1267] = 932;   M6B2[1268] = 934;   M6B2[1269] = 937;   M6B2[1270] = 939;   M6B2[1271] = 941;
    M6B2[1272] = 943;   M6B2[1273] = 945;   M6B2[1274] = 948;   M6B2[1275] = 950;   M6B2[1276] = 952;   M6B2[1277] = 954;   M6B2[1278] = 956;   M6B2[1279] = 958;
    M6B2[1280] = 896;   M6B2[1281] = 895;   M6B2[1282] = 894;   M6B2[1283] = 893;   M6B2[1284] = 892;   M6B2[1285] = 891;   M6B2[1286] = 890;   M6B2[1287] = 888;
    M6B2[1288] = 887;   M6B2[1289] = 886;   M6B2[1290] = 885;   M6B2[1291] = 884;   M6B2[1292] = 882;   M6B2[1293] = 881;   M6B2[1294] = 879;   M6B2[1295] = 878;
    M6B2[1296] = 877;   M6B2[1297] = 875;   M6B2[1298] = 874;   M6B2[1299] = 872;   M6B2[1300] = 870;   M6B2[1301] = 869;   M6B2[1302] = 867;   M6B2[1303] = 865;
    M6B2[1304] = 863;   M6B2[1305] = 862;   M6B2[1306] = 860;   M6B2[1307] = 858;   M6B2[1308] = 856;   M6B2[1309] = 853;   M6B2[1310] = 851;   M6B2[1311] = 849;
    M6B2[1312] = 847;   M6B2[1313] = 844;   M6B2[1314] = 842;   M6B2[1315] = 839;   M6B2[1316] = 836;   M6B2[1317] = 833;   M6B2[1318] = 830;   M6B2[1319] = 827;
    M6B2[1320] = 824;   M6B2[1321] = 820;   M6B2[1322] = 817;   M6B2[1323] = 813;   M6B2[1324] = 809;   M6B2[1325] = 805;   M6B2[1326] = 800;   M6B2[1327] = 795;
    M6B2[1328] = 790;   M6B2[1329] = 785;   M6B2[1330] = 779;   M6B2[1331] = 773;   M6B2[1332] = 766;   M6B2[1333] = 758;   M6B2[1334] = 750;   M6B2[1335] = 741;
    M6B2[1336] = 730;   M6B2[1337] = 718;   M6B2[1338] = 705;   M6B2[1339] = 688;   M6B2[1340] = 668;   M6B2[1341] = 642;   M6B2[1342] = 605;   M6B2[1343] = 542;
    M6B2[1344] = 896;   M6B2[1345] = 898;   M6B2[1346] = 900;   M6B2[1347] = 902;   M6B2[1348] = 904;   M6B2[1349] = 906;   M6B2[1350] = 908;   M6B2[1351] = 910;
    M6B2[1352] = 911;   M6B2[1353] = 913;   M6B2[1354] = 915;   M6B2[1355] = 917;   M6B2[1356] = 919;   M6B2[1357] = 920;   M6B2[1358] = 922;   M6B2[1359] = 924;
    M6B2[1360] = 926;   M6B2[1361] = 927;   M6B2[1362] = 929;   M6B2[1363] = 931;   M6B2[1364] = 932;   M6B2[1365] = 934;   M6B2[1366] = 936;   M6B2[1367] = 937;
    M6B2[1368] = 939;   M6B2[1369] = 941;   M6B2[1370] = 942;   M6B2[1371] = 944;   M6B2[1372] = 945;   M6B2[1373] = 947;   M6B2[1374] = 949;   M6B2[1375] = 950;
    M6B2[1376] = 952;   M6B2[1377] = 953;   M6B2[1378] = 955;   M6B2[1379] = 956;   M6B2[1380] = 958;   M6B2[1381] = 959;   M6B2[1382] = 961;   M6B2[1383] = 962;
    M6B2[1384] = 964;   M6B2[1385] = 965;   M6B2[1386] = 967;   M6B2[1387] = 968;   M6B2[1388] = 970;   M6B2[1389] = 971;   M6B2[1390] = 973;   M6B2[1391] = 974;
    M6B2[1392] = 975;   M6B2[1393] = 977;   M6B2[1394] = 978;   M6B2[1395] = 980;   M6B2[1396] = 981;   M6B2[1397] = 982;   M6B2[1398] = 984;   M6B2[1399] = 985;
    M6B2[1400] = 987;   M6B2[1401] = 988;   M6B2[1402] = 989;   M6B2[1403] = 991;   M6B2[1404] = 992;   M6B2[1405] = 993;   M6B2[1406] = 995;   M6B2[1407] = 996;
    M6B2[1408] = 933;   M6B2[1409] = 933;   M6B2[1410] = 933;   M6B2[1411] = 932;   M6B2[1412] = 932;   M6B2[1413] = 932;   M6B2[1414] = 931;   M6B2[1415] = 931;
    M6B2[1416] = 931;   M6B2[1417] = 930;   M6B2[1418] = 930;   M6B2[1419] = 929;   M6B2[1420] = 929;   M6B2[1421] = 929;   M6B2[1422] = 928;   M6B2[1423] = 928;
    M6B2[1424] = 927;   M6B2[1425] = 927;   M6B2[1426] = 927;   M6B2[1427] = 926;   M6B2[1428] = 926;   M6B2[1429] = 925;   M6B2[1430] = 925;   M6B2[1431] = 924;
    M6B2[1432] = 924;   M6B2[1433] = 923;   M6B2[1434] = 923;   M6B2[1435] = 922;   M6B2[1436] = 922;   M6B2[1437] = 921;   M6B2[1438] = 921;   M6B2[1439] = 920;
    M6B2[1440] = 920;   M6B2[1441] = 919;   M6B2[1442] = 919;   M6B2[1443] = 918;   M6B2[1444] = 917;   M6B2[1445] = 917;   M6B2[1446] = 916;   M6B2[1447] = 916;
    M6B2[1448] = 915;   M6B2[1449] = 914;   M6B2[1450] = 914;   M6B2[1451] = 913;   M6B2[1452] = 912;   M6B2[1453] = 912;   M6B2[1454] = 911;   M6B2[1455] = 910;
    M6B2[1456] = 910;   M6B2[1457] = 909;   M6B2[1458] = 908;   M6B2[1459] = 907;   M6B2[1460] = 907;   M6B2[1461] = 906;   M6B2[1462] = 905;   M6B2[1463] = 904;
    M6B2[1464] = 903;   M6B2[1465] = 903;   M6B2[1466] = 902;   M6B2[1467] = 901;   M6B2[1468] = 900;   M6B2[1469] = 899;   M6B2[1470] = 898;   M6B2[1471] = 897;
    M6B2[1472] = 933;   M6B2[1473] = 935;   M6B2[1474] = 936;   M6B2[1475] = 937;   M6B2[1476] = 939;   M6B2[1477] = 940;   M6B2[1478] = 941;   M6B2[1479] = 943;
    M6B2[1480] = 944;   M6B2[1481] = 945;   M6B2[1482] = 947;   M6B2[1483] = 948;   M6B2[1484] = 949;   M6B2[1485] = 950;   M6B2[1486] = 952;   M6B2[1487] = 953;
    M6B2[1488] = 954;   M6B2[1489] = 955;   M6B2[1490] = 957;   M6B2[1491] = 958;   M6B2[1492] = 959;   M6B2[1493] = 960;   M6B2[1494] = 962;   M6B2[1495] = 963;
    M6B2[1496] = 964;   M6B2[1497] = 965;   M6B2[1498] = 967;   M6B2[1499] = 968;   M6B2[1500] = 969;   M6B2[1501] = 970;   M6B2[1502] = 972;   M6B2[1503] = 973;
    M6B2[1504] = 974;   M6B2[1505] = 975;   M6B2[1506] = 976;   M6B2[1507] = 978;   M6B2[1508] = 979;   M6B2[1509] = 980;   M6B2[1510] = 981;   M6B2[1511] = 982;
    M6B2[1512] = 984;   M6B2[1513] = 985;   M6B2[1514] = 986;   M6B2[1515] = 987;   M6B2[1516] = 988;   M6B2[1517] = 990;   M6B2[1518] = 991;   M6B2[1519] = 992;
    M6B2[1520] = 993;   M6B2[1521] = 994;   M6B2[1522] = 995;   M6B2[1523] = 997;   M6B2[1524] = 998;   M6B2[1525] = 999;   M6B2[1526] = 1000;   M6B2[1527] = 1001;
    M6B2[1528] = 1002;   M6B2[1529] = 1004;   M6B2[1530] = 1005;   M6B2[1531] = 1006;   M6B2[1532] = 1007;   M6B2[1533] = 1008;   M6B2[1534] = 1009;   M6B2[1535] = 1011;
    M6B2[1536] = 948;   M6B2[1537] = 948;   M6B2[1538] = 947;   M6B2[1539] = 947;   M6B2[1540] = 947;   M6B2[1541] = 947;   M6B2[1542] = 947;   M6B2[1543] = 947;
    M6B2[1544] = 946;   M6B2[1545] = 946;   M6B2[1546] = 946;   M6B2[1547] = 946;   M6B2[1548] = 946;   M6B2[1549] = 946;   M6B2[1550] = 945;   M6B2[1551] = 945;
    M6B2[1552] = 945;   M6B2[1553] = 945;   M6B2[1554] = 945;   M6B2[1555] = 945;   M6B2[1556] = 944;   M6B2[1557] = 944;   M6B2[1558] = 944;   M6B2[1559] = 944;
    M6B2[1560] = 944;   M6B2[1561] = 943;   M6B2[1562] = 943;   M6B2[1563] = 943;   M6B2[1564] = 943;   M6B2[1565] = 943;   M6B2[1566] = 942;   M6B2[1567] = 942;
    M6B2[1568] = 942;   M6B2[1569] = 942;   M6B2[1570] = 942;   M6B2[1571] = 941;   M6B2[1572] = 941;   M6B2[1573] = 941;   M6B2[1574] = 941;   M6B2[1575] = 940;
    M6B2[1576] = 940;   M6B2[1577] = 940;   M6B2[1578] = 940;   M6B2[1579] = 939;   M6B2[1580] = 939;   M6B2[1581] = 939;   M6B2[1582] = 939;   M6B2[1583] = 938;
    M6B2[1584] = 938;   M6B2[1585] = 938;   M6B2[1586] = 938;   M6B2[1587] = 937;   M6B2[1588] = 937;   M6B2[1589] = 937;   M6B2[1590] = 937;   M6B2[1591] = 936;
    M6B2[1592] = 936;   M6B2[1593] = 936;   M6B2[1594] = 935;   M6B2[1595] = 935;   M6B2[1596] = 935;   M6B2[1597] = 934;   M6B2[1598] = 934;   M6B2[1599] = 934;
    M6B2[1600] = 948;   M6B2[1601] = 949;   M6B2[1602] = 950;   M6B2[1603] = 951;   M6B2[1604] = 952;   M6B2[1605] = 953;   M6B2[1606] = 954;   M6B2[1607] = 956;
    M6B2[1608] = 957;   M6B2[1609] = 958;   M6B2[1610] = 959;   M6B2[1611] = 960;   M6B2[1612] = 961;   M6B2[1613] = 962;   M6B2[1614] = 964;   M6B2[1615] = 965;
    M6B2[1616] = 966;   M6B2[1617] = 967;   M6B2[1618] = 968;   M6B2[1619] = 969;   M6B2[1620] = 970;   M6B2[1621] = 971;   M6B2[1622] = 972;   M6B2[1623] = 974;
    M6B2[1624] = 975;   M6B2[1625] = 976;   M6B2[1626] = 977;   M6B2[1627] = 978;   M6B2[1628] = 979;   M6B2[1629] = 980;   M6B2[1630] = 981;   M6B2[1631] = 982;
    M6B2[1632] = 983;   M6B2[1633] = 985;   M6B2[1634] = 986;   M6B2[1635] = 987;   M6B2[1636] = 988;   M6B2[1637] = 989;   M6B2[1638] = 990;   M6B2[1639] = 991;
    M6B2[1640] = 992;   M6B2[1641] = 993;   M6B2[1642] = 994;   M6B2[1643] = 995;   M6B2[1644] = 997;   M6B2[1645] = 998;   M6B2[1646] = 999;   M6B2[1647] = 1000;
    M6B2[1648] = 1001;   M6B2[1649] = 1002;   M6B2[1650] = 1003;   M6B2[1651] = 1004;   M6B2[1652] = 1005;   M6B2[1653] = 1006;   M6B2[1654] = 1007;   M6B2[1655] = 1008;
    M6B2[1656] = 1009;   M6B2[1657] = 1011;   M6B2[1658] = 1012;   M6B2[1659] = 1013;   M6B2[1660] = 1014;   M6B2[1661] = 1015;   M6B2[1662] = 1016;   M6B2[1663] = 1017;
    M6B2[1664] = 954;   M6B2[1665] = 954;   M6B2[1666] = 954;   M6B2[1667] = 954;   M6B2[1668] = 954;   M6B2[1669] = 954;   M6B2[1670] = 954;   M6B2[1671] = 954;
    M6B2[1672] = 953;   M6B2[1673] = 953;   M6B2[1674] = 953;   M6B2[1675] = 953;   M6B2[1676] = 953;   M6B2[1677] = 953;   M6B2[1678] = 953;   M6B2[1679] = 953;
    M6B2[1680] = 953;   M6B2[1681] = 953;   M6B2[1682] = 953;   M6B2[1683] = 953;   M6B2[1684] = 953;   M6B2[1685] = 952;   M6B2[1686] = 952;   M6B2[1687] = 952;
    M6B2[1688] = 952;   M6B2[1689] = 952;   M6B2[1690] = 952;   M6B2[1691] = 952;   M6B2[1692] = 952;   M6B2[1693] = 952;   M6B2[1694] = 952;   M6B2[1695] = 952;
    M6B2[1696] = 951;   M6B2[1697] = 951;   M6B2[1698] = 951;   M6B2[1699] = 951;   M6B2[1700] = 951;   M6B2[1701] = 951;   M6B2[1702] = 951;   M6B2[1703] = 951;
    M6B2[1704] = 951;   M6B2[1705] = 951;   M6B2[1706] = 950;   M6B2[1707] = 950;   M6B2[1708] = 950;   M6B2[1709] = 950;   M6B2[1710] = 950;   M6B2[1711] = 950;
    M6B2[1712] = 950;   M6B2[1713] = 950;   M6B2[1714] = 950;   M6B2[1715] = 949;   M6B2[1716] = 949;   M6B2[1717] = 949;   M6B2[1718] = 949;   M6B2[1719] = 949;
    M6B2[1720] = 949;   M6B2[1721] = 949;   M6B2[1722] = 948;   M6B2[1723] = 948;   M6B2[1724] = 948;   M6B2[1725] = 948;   M6B2[1726] = 948;   M6B2[1727] = 948;
    M6B2[1728] = 954;   M6B2[1729] = 955;   M6B2[1730] = 956;   M6B2[1731] = 957;   M6B2[1732] = 958;   M6B2[1733] = 959;   M6B2[1734] = 960;   M6B2[1735] = 961;
    M6B2[1736] = 963;   M6B2[1737] = 964;   M6B2[1738] = 965;   M6B2[1739] = 966;   M6B2[1740] = 967;   M6B2[1741] = 968;   M6B2[1742] = 969;   M6B2[1743] = 970;
    M6B2[1744] = 971;   M6B2[1745] = 972;   M6B2[1746] = 973;   M6B2[1747] = 974;   M6B2[1748] = 975;   M6B2[1749] = 976;   M6B2[1750] = 977;   M6B2[1751] = 978;
    M6B2[1752] = 979;   M6B2[1753] = 980;   M6B2[1754] = 982;   M6B2[1755] = 983;   M6B2[1756] = 984;   M6B2[1757] = 985;   M6B2[1758] = 986;   M6B2[1759] = 987;
    M6B2[1760] = 988;   M6B2[1761] = 989;   M6B2[1762] = 990;   M6B2[1763] = 991;   M6B2[1764] = 992;   M6B2[1765] = 993;   M6B2[1766] = 994;   M6B2[1767] = 995;
    M6B2[1768] = 996;   M6B2[1769] = 997;   M6B2[1770] = 998;   M6B2[1771] = 999;   M6B2[1772] = 1000;   M6B2[1773] = 1001;   M6B2[1774] = 1002;   M6B2[1775] = 1003;
    M6B2[1776] = 1005;   M6B2[1777] = 1006;   M6B2[1778] = 1007;   M6B2[1779] = 1008;   M6B2[1780] = 1009;   M6B2[1781] = 1010;   M6B2[1782] = 1011;   M6B2[1783] = 1012;
    M6B2[1784] = 1013;   M6B2[1785] = 1014;   M6B2[1786] = 1015;   M6B2[1787] = 1016;   M6B2[1788] = 1017;   M6B2[1789] = 1018;   M6B2[1790] = 1019;   M6B2[1791] = 1020;
    M6B2[1792] = 957;   M6B2[1793] = 957;   M6B2[1794] = 957;   M6B2[1795] = 957;   M6B2[1796] = 957;   M6B2[1797] = 957;   M6B2[1798] = 957;   M6B2[1799] = 957;
    M6B2[1800] = 957;   M6B2[1801] = 957;   M6B2[1802] = 957;   M6B2[1803] = 957;   M6B2[1804] = 957;   M6B2[1805] = 957;   M6B2[1806] = 957;   M6B2[1807] = 957;
    M6B2[1808] = 957;   M6B2[1809] = 956;   M6B2[1810] = 956;   M6B2[1811] = 956;   M6B2[1812] = 956;   M6B2[1813] = 956;   M6B2[1814] = 956;   M6B2[1815] = 956;
    M6B2[1816] = 956;   M6B2[1817] = 956;   M6B2[1818] = 956;   M6B2[1819] = 956;   M6B2[1820] = 956;   M6B2[1821] = 956;   M6B2[1822] = 956;   M6B2[1823] = 956;
    M6B2[1824] = 956;   M6B2[1825] = 956;   M6B2[1826] = 956;   M6B2[1827] = 956;   M6B2[1828] = 956;   M6B2[1829] = 956;   M6B2[1830] = 956;   M6B2[1831] = 955;
    M6B2[1832] = 955;   M6B2[1833] = 955;   M6B2[1834] = 955;   M6B2[1835] = 955;   M6B2[1836] = 955;   M6B2[1837] = 955;   M6B2[1838] = 955;   M6B2[1839] = 955;
    M6B2[1840] = 955;   M6B2[1841] = 955;   M6B2[1842] = 955;   M6B2[1843] = 955;   M6B2[1844] = 955;   M6B2[1845] = 955;   M6B2[1846] = 955;   M6B2[1847] = 955;
    M6B2[1848] = 955;   M6B2[1849] = 954;   M6B2[1850] = 954;   M6B2[1851] = 954;   M6B2[1852] = 954;   M6B2[1853] = 954;   M6B2[1854] = 954;   M6B2[1855] = 954;
    M6B2[1856] = 957;   M6B2[1857] = 958;   M6B2[1858] = 959;   M6B2[1859] = 960;   M6B2[1860] = 961;   M6B2[1861] = 962;   M6B2[1862] = 963;   M6B2[1863] = 964;
    M6B2[1864] = 965;   M6B2[1865] = 966;   M6B2[1866] = 967;   M6B2[1867] = 968;   M6B2[1868] = 969;   M6B2[1869] = 970;   M6B2[1870] = 971;   M6B2[1871] = 973;
    M6B2[1872] = 974;   M6B2[1873] = 975;   M6B2[1874] = 976;   M6B2[1875] = 977;   M6B2[1876] = 978;   M6B2[1877] = 979;   M6B2[1878] = 980;   M6B2[1879] = 981;
    M6B2[1880] = 982;   M6B2[1881] = 983;   M6B2[1882] = 984;   M6B2[1883] = 985;   M6B2[1884] = 986;   M6B2[1885] = 987;   M6B2[1886] = 988;   M6B2[1887] = 989;
    M6B2[1888] = 990;   M6B2[1889] = 991;   M6B2[1890] = 992;   M6B2[1891] = 993;   M6B2[1892] = 994;   M6B2[1893] = 995;   M6B2[1894] = 996;   M6B2[1895] = 997;
    M6B2[1896] = 998;   M6B2[1897] = 999;   M6B2[1898] = 1000;   M6B2[1899] = 1001;   M6B2[1900] = 1002;   M6B2[1901] = 1003;   M6B2[1902] = 1004;   M6B2[1903] = 1005;
    M6B2[1904] = 1006;   M6B2[1905] = 1007;   M6B2[1906] = 1008;   M6B2[1907] = 1009;   M6B2[1908] = 1010;   M6B2[1909] = 1011;   M6B2[1910] = 1012;   M6B2[1911] = 1013;
    M6B2[1912] = 1014;   M6B2[1913] = 1015;   M6B2[1914] = 1016;   M6B2[1915] = 1017;   M6B2[1916] = 1018;   M6B2[1917] = 1019;   M6B2[1918] = 1021;   M6B2[1919] = 1022;
    M6B2[1920] = 959;   M6B2[1921] = 959;   M6B2[1922] = 959;   M6B2[1923] = 958;   M6B2[1924] = 958;   M6B2[1925] = 958;   M6B2[1926] = 958;   M6B2[1927] = 958;
    M6B2[1928] = 958;   M6B2[1929] = 958;   M6B2[1930] = 958;   M6B2[1931] = 958;   M6B2[1932] = 958;   M6B2[1933] = 958;   M6B2[1934] = 958;   M6B2[1935] = 958;
    M6B2[1936] = 958;   M6B2[1937] = 958;   M6B2[1938] = 958;   M6B2[1939] = 958;   M6B2[1940] = 958;   M6B2[1941] = 958;   M6B2[1942] = 958;   M6B2[1943] = 958;
    M6B2[1944] = 958;   M6B2[1945] = 958;   M6B2[1946] = 958;   M6B2[1947] = 958;   M6B2[1948] = 958;   M6B2[1949] = 958;   M6B2[1950] = 958;   M6B2[1951] = 958;
    M6B2[1952] = 958;   M6B2[1953] = 958;   M6B2[1954] = 958;   M6B2[1955] = 958;   M6B2[1956] = 958;   M6B2[1957] = 958;   M6B2[1958] = 958;   M6B2[1959] = 958;
    M6B2[1960] = 958;   M6B2[1961] = 958;   M6B2[1962] = 958;   M6B2[1963] = 958;   M6B2[1964] = 958;   M6B2[1965] = 958;   M6B2[1966] = 958;   M6B2[1967] = 958;
    M6B2[1968] = 958;   M6B2[1969] = 958;   M6B2[1970] = 957;   M6B2[1971] = 957;   M6B2[1972] = 957;   M6B2[1973] = 957;   M6B2[1974] = 957;   M6B2[1975] = 957;
    M6B2[1976] = 957;   M6B2[1977] = 957;   M6B2[1978] = 957;   M6B2[1979] = 957;   M6B2[1980] = 957;   M6B2[1981] = 957;   M6B2[1982] = 957;   M6B2[1983] = 957;
    M6B2[1984] = 959;   M6B2[1985] = 960;   M6B2[1986] = 961;   M6B2[1987] = 962;   M6B2[1988] = 963;   M6B2[1989] = 964;   M6B2[1990] = 965;   M6B2[1991] = 966;
    M6B2[1992] = 967;   M6B2[1993] = 968;   M6B2[1994] = 969;   M6B2[1995] = 970;   M6B2[1996] = 971;   M6B2[1997] = 972;   M6B2[1998] = 973;   M6B2[1999] = 974;
    M6B2[2000] = 975;   M6B2[2001] = 976;   M6B2[2002] = 977;   M6B2[2003] = 978;   M6B2[2004] = 979;   M6B2[2005] = 980;   M6B2[2006] = 981;   M6B2[2007] = 982;
    M6B2[2008] = 983;   M6B2[2009] = 984;   M6B2[2010] = 985;   M6B2[2011] = 986;   M6B2[2012] = 987;   M6B2[2013] = 988;   M6B2[2014] = 989;   M6B2[2015] = 990;
    M6B2[2016] = 991;   M6B2[2017] = 992;   M6B2[2018] = 993;   M6B2[2019] = 994;   M6B2[2020] = 995;   M6B2[2021] = 996;   M6B2[2022] = 997;   M6B2[2023] = 998;
    M6B2[2024] = 999;   M6B2[2025] = 1000;   M6B2[2026] = 1001;   M6B2[2027] = 1002;   M6B2[2028] = 1003;   M6B2[2029] = 1004;   M6B2[2030] = 1005;   M6B2[2031] = 1006;
    M6B2[2032] = 1007;   M6B2[2033] = 1008;   M6B2[2034] = 1009;   M6B2[2035] = 1010;   M6B2[2036] = 1011;   M6B2[2037] = 1012;   M6B2[2038] = 1013;   M6B2[2039] = 1014;
    M6B2[2040] = 1015;   M6B2[2041] = 1016;   M6B2[2042] = 1017;   M6B2[2043] = 1018;   M6B2[2044] = 1019;   M6B2[2045] = 1020;   M6B2[2046] = 1021;   M6B2[2047] = 1022;
    M6B2[2048] = 959;   M6B2[2049] = 959;   M6B2[2050] = 959;   M6B2[2051] = 959;   M6B2[2052] = 959;   M6B2[2053] = 959;   M6B2[2054] = 959;   M6B2[2055] = 959;
    M6B2[2056] = 959;   M6B2[2057] = 959;   M6B2[2058] = 959;   M6B2[2059] = 959;   M6B2[2060] = 959;   M6B2[2061] = 959;   M6B2[2062] = 959;   M6B2[2063] = 959;
    M6B2[2064] = 959;   M6B2[2065] = 959;   M6B2[2066] = 959;   M6B2[2067] = 959;   M6B2[2068] = 959;   M6B2[2069] = 959;   M6B2[2070] = 959;   M6B2[2071] = 959;
    M6B2[2072] = 959;   M6B2[2073] = 959;   M6B2[2074] = 959;   M6B2[2075] = 959;   M6B2[2076] = 959;   M6B2[2077] = 959;   M6B2[2078] = 959;   M6B2[2079] = 959;
    M6B2[2080] = 959;   M6B2[2081] = 959;   M6B2[2082] = 959;   M6B2[2083] = 959;   M6B2[2084] = 959;   M6B2[2085] = 959;   M6B2[2086] = 959;   M6B2[2087] = 959;
    M6B2[2088] = 959;   M6B2[2089] = 959;   M6B2[2090] = 959;   M6B2[2091] = 959;   M6B2[2092] = 959;   M6B2[2093] = 959;   M6B2[2094] = 959;   M6B2[2095] = 959;
    M6B2[2096] = 959;   M6B2[2097] = 959;   M6B2[2098] = 959;   M6B2[2099] = 959;   M6B2[2100] = 959;   M6B2[2101] = 959;   M6B2[2102] = 959;   M6B2[2103] = 959;
    M6B2[2104] = 959;   M6B2[2105] = 959;   M6B2[2106] = 959;   M6B2[2107] = 959;   M6B2[2108] = 959;   M6B2[2109] = 959;   M6B2[2110] = 959;   M6B2[2111] = 959;
    M6B2[2112] = 959;   M6B2[2113] = 960;   M6B2[2114] = 961;   M6B2[2115] = 962;   M6B2[2116] = 963;   M6B2[2117] = 964;   M6B2[2118] = 965;   M6B2[2119] = 966;
    M6B2[2120] = 967;   M6B2[2121] = 968;   M6B2[2122] = 969;   M6B2[2123] = 970;   M6B2[2124] = 971;   M6B2[2125] = 972;   M6B2[2126] = 973;   M6B2[2127] = 974;
    M6B2[2128] = 975;   M6B2[2129] = 976;   M6B2[2130] = 977;   M6B2[2131] = 978;   M6B2[2132] = 979;   M6B2[2133] = 980;   M6B2[2134] = 981;   M6B2[2135] = 982;
    M6B2[2136] = 983;   M6B2[2137] = 984;   M6B2[2138] = 985;   M6B2[2139] = 986;   M6B2[2140] = 987;   M6B2[2141] = 988;   M6B2[2142] = 989;   M6B2[2143] = 990;
    M6B2[2144] = 991;   M6B2[2145] = 992;   M6B2[2146] = 993;   M6B2[2147] = 995;   M6B2[2148] = 996;   M6B2[2149] = 997;   M6B2[2150] = 998;   M6B2[2151] = 999;
    M6B2[2152] = 1000;   M6B2[2153] = 1001;   M6B2[2154] = 1002;   M6B2[2155] = 1003;   M6B2[2156] = 1004;   M6B2[2157] = 1005;   M6B2[2158] = 1006;   M6B2[2159] = 1007;
    M6B2[2160] = 1008;   M6B2[2161] = 1009;   M6B2[2162] = 1010;   M6B2[2163] = 1011;   M6B2[2164] = 1012;   M6B2[2165] = 1013;   M6B2[2166] = 1014;   M6B2[2167] = 1015;
    M6B2[2168] = 1016;   M6B2[2169] = 1017;   M6B2[2170] = 1018;   M6B2[2171] = 1019;   M6B2[2172] = 1020;   M6B2[2173] = 1021;   M6B2[2174] = 1022;   M6B2[2175] = 1023;
    M6B2[2176] = 960;   M6B2[2177] = 960;   M6B2[2178] = 960;   M6B2[2179] = 960;   M6B2[2180] = 960;   M6B2[2181] = 960;   M6B2[2182] = 960;   M6B2[2183] = 960;
    M6B2[2184] = 960;   M6B2[2185] = 960;   M6B2[2186] = 960;   M6B2[2187] = 960;   M6B2[2188] = 960;   M6B2[2189] = 960;   M6B2[2190] = 960;   M6B2[2191] = 960;
    M6B2[2192] = 960;   M6B2[2193] = 960;   M6B2[2194] = 960;   M6B2[2195] = 960;   M6B2[2196] = 960;   M6B2[2197] = 960;   M6B2[2198] = 960;   M6B2[2199] = 960;
    M6B2[2200] = 960;   M6B2[2201] = 960;   M6B2[2202] = 960;   M6B2[2203] = 960;   M6B2[2204] = 960;   M6B2[2205] = 960;   M6B2[2206] = 959;   M6B2[2207] = 959;
    M6B2[2208] = 959;   M6B2[2209] = 959;   M6B2[2210] = 959;   M6B2[2211] = 959;   M6B2[2212] = 959;   M6B2[2213] = 959;   M6B2[2214] = 959;   M6B2[2215] = 959;
    M6B2[2216] = 959;   M6B2[2217] = 959;   M6B2[2218] = 959;   M6B2[2219] = 959;   M6B2[2220] = 959;   M6B2[2221] = 959;   M6B2[2222] = 959;   M6B2[2223] = 959;
    M6B2[2224] = 959;   M6B2[2225] = 959;   M6B2[2226] = 959;   M6B2[2227] = 959;   M6B2[2228] = 959;   M6B2[2229] = 959;   M6B2[2230] = 959;   M6B2[2231] = 959;
    M6B2[2232] = 959;   M6B2[2233] = 959;   M6B2[2234] = 959;   M6B2[2235] = 959;   M6B2[2236] = 959;   M6B2[2237] = 959;   M6B2[2238] = 959;   M6B2[2239] = 959;
    M6B2[2240] = 960;   M6B2[2241] = 961;   M6B2[2242] = 962;   M6B2[2243] = 963;   M6B2[2244] = 964;   M6B2[2245] = 965;   M6B2[2246] = 966;   M6B2[2247] = 967;
    M6B2[2248] = 968;   M6B2[2249] = 969;   M6B2[2250] = 970;   M6B2[2251] = 971;   M6B2[2252] = 972;   M6B2[2253] = 973;   M6B2[2254] = 974;   M6B2[2255] = 975;
    M6B2[2256] = 976;   M6B2[2257] = 977;   M6B2[2258] = 978;   M6B2[2259] = 979;   M6B2[2260] = 980;   M6B2[2261] = 981;   M6B2[2262] = 982;   M6B2[2263] = 983;
    M6B2[2264] = 984;   M6B2[2265] = 985;   M6B2[2266] = 986;   M6B2[2267] = 987;   M6B2[2268] = 988;   M6B2[2269] = 989;   M6B2[2270] = 990;   M6B2[2271] = 991;
    M6B2[2272] = 992;   M6B2[2273] = 993;   M6B2[2274] = 994;   M6B2[2275] = 995;   M6B2[2276] = 996;   M6B2[2277] = 997;   M6B2[2278] = 998;   M6B2[2279] = 999;
    M6B2[2280] = 1000;   M6B2[2281] = 1001;   M6B2[2282] = 1002;   M6B2[2283] = 1003;   M6B2[2284] = 1004;   M6B2[2285] = 1005;   M6B2[2286] = 1006;   M6B2[2287] = 1007;
    M6B2[2288] = 1008;   M6B2[2289] = 1009;   M6B2[2290] = 1010;   M6B2[2291] = 1011;   M6B2[2292] = 1012;   M6B2[2293] = 1013;   M6B2[2294] = 1014;   M6B2[2295] = 1015;
    M6B2[2296] = 1016;   M6B2[2297] = 1017;   M6B2[2298] = 1018;   M6B2[2299] = 1019;   M6B2[2300] = 1020;   M6B2[2301] = 1021;   M6B2[2302] = 1022;   M6B2[2303] = 1023;
end

// 根据最大位数选择对应的数组并进行查找
always @(*) begin
    case(max_bit)
        5'd1: begin
            // for (j = 0; j < 4; j = j + 1) begin
            //     for (i = 0; i < 8; i = i + 1) begin
            //         lookup_result_0[j][i] = M1B2[addra[j][i]];
            //     end
            // end
        end
        5'd2: begin
            // for (j = 0; j < 4; j = j + 1) begin
            //     for (i = 0; i < 8; i = i + 1) begin
            //         lookup_result_0[j][i] = M2B2[addra[j][i]];
            //     end
            // end
        end
        5'd3: begin
            // for (j = 0; j < 4; j = j + 1) begin
            //     for (i = 0; i < 8; i = i + 1) begin
            //         lookup_result_0[j][i] = M3B2[addra[j][i]];
            //     end
            // end
        end
        5'd4: begin
            // for (j = 0; j < 4; j = j + 1) begin
            //     for (i = 0; i < 8; i = i + 1) begin
            //         lookup_result_0[j][i] = M4B2[addra[j][i]];
            //     end
            // end
        end
        5'd5: begin            
            // for (j = 0; j < 4; j = j + 1) begin
            //     for (i = 0; i < 8; i = i + 1) begin
            //         lookup_result_0[j][i] = M5B2[addra[j][i]];
            //     end
            // end
        end
        5'd6: begin            
            for (j = 0; j < 4; j = j + 1) begin
                for (i = 0; i < 8; i = i + 1) begin
                    lookup_result_0[j][i] = M6B2[addra[j][i]];
                end
            end
        end
        default: begin

        end
    endcase
end
// 将查找结果连接到输出
assign result_bin = lookup_result_0;
endmodule
